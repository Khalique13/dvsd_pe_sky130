magic
tech sky130A
magscale 1 2
timestamp 1633581810
<< nwell >>
rect 1066 116677 178886 117243
rect 1066 115589 178886 116155
rect 1066 114501 178886 115067
rect 1066 113413 178886 113979
rect 1066 112325 178886 112891
rect 1066 111237 178886 111803
rect 1066 110149 178886 110715
rect 1066 109061 178886 109627
rect 1066 107973 178886 108539
rect 1066 106885 178886 107451
rect 1066 105797 178886 106363
rect 1066 104709 178886 105275
rect 1066 103621 178886 104187
rect 1066 102533 178886 103099
rect 1066 101445 178886 102011
rect 1066 100357 178886 100923
rect 1066 99269 178886 99835
rect 1066 98181 178886 98747
rect 1066 97093 178886 97659
rect 1066 96005 178886 96571
rect 1066 94917 178886 95483
rect 1066 93829 178886 94395
rect 1066 92741 178886 93307
rect 1066 91653 178886 92219
rect 1066 90565 178886 91131
rect 1066 89477 178886 90043
rect 1066 88389 178886 88955
rect 1066 87301 178886 87867
rect 1066 86213 178886 86779
rect 1066 85125 178886 85691
rect 1066 84037 178886 84603
rect 1066 82949 178886 83515
rect 1066 81861 178886 82427
rect 1066 80773 178886 81339
rect 1066 79685 178886 80251
rect 1066 78597 178886 79163
rect 1066 77509 178886 78075
rect 1066 76421 178886 76987
rect 1066 75333 178886 75899
rect 1066 74245 178886 74811
rect 1066 73157 178886 73723
rect 1066 72069 178886 72635
rect 1066 70981 178886 71547
rect 1066 69893 178886 70459
rect 1066 68805 178886 69371
rect 1066 67717 178886 68283
rect 1066 66629 178886 67195
rect 1066 65541 178886 66107
rect 1066 64453 178886 65019
rect 1066 63365 178886 63931
rect 1066 62277 178886 62843
rect 1066 61189 178886 61755
rect 1066 60101 178886 60667
rect 1066 59013 178886 59579
rect 1066 57925 178886 58491
rect 1066 56837 178886 57403
rect 1066 55749 178886 56315
rect 1066 54661 178886 55227
rect 1066 53573 178886 54139
rect 1066 52485 178886 53051
rect 1066 51397 178886 51963
rect 1066 50309 178886 50875
rect 1066 49221 178886 49787
rect 1066 48133 178886 48699
rect 1066 47045 178886 47611
rect 1066 45957 178886 46523
rect 1066 44869 178886 45435
rect 1066 43781 178886 44347
rect 1066 42693 178886 43259
rect 1066 41605 178886 42171
rect 1066 40517 178886 41083
rect 1066 39429 178886 39995
rect 1066 38341 178886 38907
rect 1066 37253 178886 37819
rect 1066 36165 178886 36731
rect 1066 35077 178886 35643
rect 1066 33989 178886 34555
rect 1066 32901 178886 33467
rect 1066 31813 178886 32379
rect 1066 30725 178886 31291
rect 1066 29637 178886 30203
rect 1066 28549 178886 29115
rect 1066 27461 178886 28027
rect 1066 26373 178886 26939
rect 1066 25285 178886 25851
rect 1066 24197 178886 24763
rect 1066 23109 178886 23675
rect 1066 22021 178886 22587
rect 1066 20933 178886 21499
rect 1066 19845 178886 20411
rect 1066 18757 178886 19323
rect 1066 17669 178886 18235
rect 1066 16581 178886 17147
rect 1066 15493 178886 16059
rect 1066 14405 178886 14971
rect 1066 13317 178886 13883
rect 1066 12229 178886 12795
rect 1066 11141 178886 11707
rect 1066 10053 178886 10619
rect 1066 8965 178886 9531
rect 1066 7877 178886 8443
rect 1066 6789 178886 7355
rect 1066 5701 178886 6267
rect 1066 4613 178886 5179
rect 1066 3525 178886 4091
rect 1066 2437 178886 3003
<< obsli1 >>
rect 1104 2159 178848 117521
<< obsm1 >>
rect 1104 2128 178848 117552
<< metal2 >>
rect 7470 119200 7526 120000
rect 22466 119200 22522 120000
rect 37462 119200 37518 120000
rect 52458 119200 52514 120000
rect 67454 119200 67510 120000
rect 82450 119200 82506 120000
rect 97446 119200 97502 120000
rect 112442 119200 112498 120000
rect 127438 119200 127494 120000
rect 142434 119200 142490 120000
rect 157430 119200 157486 120000
rect 172426 119200 172482 120000
rect 45006 0 45062 800
rect 134982 0 135038 800
<< obsm2 >>
rect 4214 119144 7414 119200
rect 7582 119144 22410 119200
rect 22578 119144 37406 119200
rect 37574 119144 52402 119200
rect 52570 119144 67398 119200
rect 67566 119144 82394 119200
rect 82562 119144 97390 119200
rect 97558 119144 112386 119200
rect 112554 119144 127382 119200
rect 127550 119144 142378 119200
rect 142546 119144 157374 119200
rect 157542 119144 172370 119200
rect 172538 119144 173482 119200
rect 4214 856 173482 119144
rect 4214 800 44950 856
rect 45118 800 134926 856
rect 135094 800 173482 856
<< obsm3 >>
rect 4208 2143 173488 117537
<< metal4 >>
rect 4208 2128 4528 117552
rect 19568 2128 19888 117552
rect 34928 2128 35248 117552
rect 50288 2128 50608 117552
rect 65648 2128 65968 117552
rect 81008 2128 81328 117552
rect 96368 2128 96688 117552
rect 111728 2128 112048 117552
rect 127088 2128 127408 117552
rect 142448 2128 142768 117552
rect 157808 2128 158128 117552
rect 173168 2128 173488 117552
<< labels >>
rlabel metal2 s 7470 119200 7526 120000 6 io_en
port 1 nsew signal input
rlabel metal2 s 22466 119200 22522 120000 6 io_in[0]
port 2 nsew signal input
rlabel metal2 s 52458 119200 52514 120000 6 io_in[1]
port 3 nsew signal input
rlabel metal2 s 82450 119200 82506 120000 6 io_in[2]
port 4 nsew signal input
rlabel metal2 s 112442 119200 112498 120000 6 io_in[3]
port 5 nsew signal input
rlabel metal2 s 127438 119200 127494 120000 6 io_in[4]
port 6 nsew signal input
rlabel metal2 s 142434 119200 142490 120000 6 io_in[5]
port 7 nsew signal input
rlabel metal2 s 157430 119200 157486 120000 6 io_in[6]
port 8 nsew signal input
rlabel metal2 s 172426 119200 172482 120000 6 io_in[7]
port 9 nsew signal input
rlabel metal2 s 37462 119200 37518 120000 6 io_out[0]
port 10 nsew signal output
rlabel metal2 s 67454 119200 67510 120000 6 io_out[1]
port 11 nsew signal output
rlabel metal2 s 97446 119200 97502 120000 6 io_out[2]
port 12 nsew signal output
rlabel metal4 s 4208 2128 4528 117552 6 vccd1
port 13 nsew power input
rlabel metal4 s 34928 2128 35248 117552 6 vccd1
port 13 nsew power input
rlabel metal4 s 65648 2128 65968 117552 6 vccd1
port 13 nsew power input
rlabel metal4 s 96368 2128 96688 117552 6 vccd1
port 13 nsew power input
rlabel metal4 s 127088 2128 127408 117552 6 vccd1
port 13 nsew power input
rlabel metal4 s 157808 2128 158128 117552 6 vccd1
port 13 nsew power input
rlabel metal4 s 19568 2128 19888 117552 6 vssd1
port 14 nsew ground input
rlabel metal4 s 50288 2128 50608 117552 6 vssd1
port 14 nsew ground input
rlabel metal4 s 81008 2128 81328 117552 6 vssd1
port 14 nsew ground input
rlabel metal4 s 111728 2128 112048 117552 6 vssd1
port 14 nsew ground input
rlabel metal4 s 142448 2128 142768 117552 6 vssd1
port 14 nsew ground input
rlabel metal4 s 173168 2128 173488 117552 6 vssd1
port 14 nsew ground input
rlabel metal2 s 45006 0 45062 800 6 wb_eno
port 15 nsew signal output
rlabel metal2 s 134982 0 135038 800 6 wb_gs
port 16 nsew signal output
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 180000 120000
string LEFview TRUE
string GDS_FILE /project/openlane/user_proj_example/runs/user_proj_example/results/magic/user_proj_example.gds
string GDS_END 5525326
string GDS_START 119578
<< end >>

