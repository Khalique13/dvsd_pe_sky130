magic
tech sky130A
magscale 1 2
timestamp 1629374141
<< locali >>
rect 5825 3519 5859 5797
rect 5917 3723 5951 8381
rect 6009 3043 6043 8449
<< viali >>
rect 1501 8585 1535 8619
rect 2145 8517 2179 8551
rect 1593 8449 1627 8483
rect 2329 8449 2363 8483
rect 3249 8449 3283 8483
rect 3985 8449 4019 8483
rect 4813 8449 4847 8483
rect 6009 8449 6043 8483
rect 5917 8381 5951 8415
rect 3157 8313 3191 8347
rect 3893 8245 3927 8279
rect 4905 8245 4939 8279
rect 1777 8041 1811 8075
rect 4261 7973 4295 8007
rect 4813 7973 4847 8007
rect 2513 7837 2547 7871
rect 2789 7837 2823 7871
rect 3985 7837 4019 7871
rect 4077 7837 4111 7871
rect 4353 7837 4387 7871
rect 4997 7837 5031 7871
rect 3801 7701 3835 7735
rect 2513 7497 2547 7531
rect 4169 7497 4203 7531
rect 1777 7361 1811 7395
rect 3249 7361 3283 7395
rect 3433 7361 3467 7395
rect 3709 7361 3743 7395
rect 4353 7361 4387 7395
rect 4813 7361 4847 7395
rect 1501 7293 1535 7327
rect 4537 7293 4571 7327
rect 3525 7225 3559 7259
rect 2973 7157 3007 7191
rect 3341 7157 3375 7191
rect 4445 7157 4479 7191
rect 2237 6953 2271 6987
rect 3985 6953 4019 6987
rect 2973 6885 3007 6919
rect 2237 6817 2271 6851
rect 2329 6817 2363 6851
rect 2881 6817 2915 6851
rect 1409 6749 1443 6783
rect 2421 6749 2455 6783
rect 3065 6749 3099 6783
rect 3157 6749 3191 6783
rect 4077 6749 4111 6783
rect 4169 6749 4203 6783
rect 4905 6749 4939 6783
rect 2053 6681 2087 6715
rect 1593 6613 1627 6647
rect 3801 6613 3835 6647
rect 4721 6613 4755 6647
rect 2887 6409 2921 6443
rect 4721 6409 4755 6443
rect 2031 6341 2065 6375
rect 2973 6341 3007 6375
rect 4077 6341 4111 6375
rect 2329 6273 2363 6307
rect 2789 6273 2823 6307
rect 3065 6273 3099 6307
rect 3801 6273 3835 6307
rect 4537 6273 4571 6307
rect 2145 6205 2179 6239
rect 2237 6205 2271 6239
rect 3893 6205 3927 6239
rect 1961 6137 1995 6171
rect 3617 6069 3651 6103
rect 4077 6069 4111 6103
rect 1685 5865 1719 5899
rect 5825 5797 5859 5831
rect 2237 5729 2271 5763
rect 3985 5729 4019 5763
rect 4353 5729 4387 5763
rect 1409 5661 1443 5695
rect 1685 5661 1719 5695
rect 2513 5661 2547 5695
rect 4077 5661 4111 5695
rect 4445 5593 4479 5627
rect 1501 5525 1535 5559
rect 3249 5525 3283 5559
rect 3801 5525 3835 5559
rect 2421 5321 2455 5355
rect 3617 5321 3651 5355
rect 1409 5253 1443 5287
rect 2605 5253 2639 5287
rect 4813 5253 4847 5287
rect 1593 5185 1627 5219
rect 1777 5185 1811 5219
rect 2789 5185 2823 5219
rect 3985 5185 4019 5219
rect 3893 5117 3927 5151
rect 4997 5049 5031 5083
rect 3801 4981 3835 5015
rect 1409 4777 1443 4811
rect 2605 4777 2639 4811
rect 3801 4777 3835 4811
rect 2973 4709 3007 4743
rect 1869 4641 1903 4675
rect 2697 4641 2731 4675
rect 4445 4641 4479 4675
rect 1685 4573 1719 4607
rect 1777 4573 1811 4607
rect 2145 4573 2179 4607
rect 2605 4573 2639 4607
rect 3926 4573 3960 4607
rect 4353 4573 4387 4607
rect 2053 4437 2087 4471
rect 3985 4437 4019 4471
rect 3525 4233 3559 4267
rect 4445 4233 4479 4267
rect 2145 4097 2179 4131
rect 2605 4097 2639 4131
rect 3709 4097 3743 4131
rect 4261 4097 4295 4131
rect 1869 4029 1903 4063
rect 2421 3961 2455 3995
rect 2237 3893 2271 3927
rect 2329 3893 2363 3927
rect 1593 3689 1627 3723
rect 2145 3689 2179 3723
rect 2329 3689 2363 3723
rect 3893 3689 3927 3723
rect 4813 3689 4847 3723
rect 2421 3553 2455 3587
rect 5917 3689 5951 3723
rect 1501 3485 1535 3519
rect 2697 3485 2731 3519
rect 3801 3485 3835 3519
rect 4997 3485 5031 3519
rect 5825 3485 5859 3519
rect 1593 3145 1627 3179
rect 2881 3145 2915 3179
rect 3617 3145 3651 3179
rect 4353 3145 4387 3179
rect 1409 3009 1443 3043
rect 2145 3009 2179 3043
rect 2329 3009 2363 3043
rect 2789 3009 2823 3043
rect 3433 3009 3467 3043
rect 4169 3009 4203 3043
rect 4813 3009 4847 3043
rect 6009 3009 6043 3043
rect 2237 2873 2271 2907
rect 4905 2805 4939 2839
rect 2881 2601 2915 2635
rect 4261 2601 4295 2635
rect 1685 2465 1719 2499
rect 1409 2397 1443 2431
rect 2697 2397 2731 2431
rect 4077 2397 4111 2431
rect 4813 2397 4847 2431
rect 4997 2329 5031 2363
<< metal1 >>
rect 1104 8730 5704 8752
rect 1104 8678 2523 8730
rect 2575 8678 2587 8730
rect 2639 8678 2651 8730
rect 2703 8678 2715 8730
rect 2767 8678 4065 8730
rect 4117 8678 4129 8730
rect 4181 8678 4193 8730
rect 4245 8678 4257 8730
rect 4309 8678 5704 8730
rect 1104 8656 5704 8678
rect 1486 8616 1492 8628
rect 1447 8588 1492 8616
rect 1486 8576 1492 8588
rect 1544 8576 1550 8628
rect 566 8508 572 8560
rect 624 8548 630 8560
rect 2133 8551 2191 8557
rect 2133 8548 2145 8551
rect 624 8520 2145 8548
rect 624 8508 630 8520
rect 2133 8517 2145 8520
rect 2179 8517 2191 8551
rect 2133 8511 2191 8517
rect 1578 8480 1584 8492
rect 1539 8452 1584 8480
rect 1578 8440 1584 8452
rect 1636 8440 1642 8492
rect 2314 8480 2320 8492
rect 2275 8452 2320 8480
rect 2314 8440 2320 8452
rect 2372 8440 2378 8492
rect 3237 8483 3295 8489
rect 3237 8449 3249 8483
rect 3283 8449 3295 8483
rect 3237 8443 3295 8449
rect 3252 8412 3280 8443
rect 3878 8440 3884 8492
rect 3936 8480 3942 8492
rect 3973 8483 4031 8489
rect 3973 8480 3985 8483
rect 3936 8452 3985 8480
rect 3936 8440 3942 8452
rect 3973 8449 3985 8452
rect 4019 8449 4031 8483
rect 3973 8443 4031 8449
rect 4801 8483 4859 8489
rect 4801 8449 4813 8483
rect 4847 8480 4859 8483
rect 5997 8483 6055 8489
rect 5997 8480 6009 8483
rect 4847 8452 6009 8480
rect 4847 8449 4859 8452
rect 4801 8443 4859 8449
rect 5997 8449 6009 8452
rect 6043 8449 6055 8483
rect 5997 8443 6055 8449
rect 4706 8412 4712 8424
rect 3252 8384 4712 8412
rect 4706 8372 4712 8384
rect 4764 8412 4770 8424
rect 5905 8415 5963 8421
rect 5905 8412 5917 8415
rect 4764 8384 5917 8412
rect 4764 8372 4770 8384
rect 5905 8381 5917 8384
rect 5951 8381 5963 8415
rect 5905 8375 5963 8381
rect 3145 8347 3203 8353
rect 3145 8313 3157 8347
rect 3191 8344 3203 8347
rect 4062 8344 4068 8356
rect 3191 8316 4068 8344
rect 3191 8313 3203 8316
rect 3145 8307 3203 8313
rect 4062 8304 4068 8316
rect 4120 8304 4126 8356
rect 3602 8236 3608 8288
rect 3660 8276 3666 8288
rect 3881 8279 3939 8285
rect 3881 8276 3893 8279
rect 3660 8248 3893 8276
rect 3660 8236 3666 8248
rect 3881 8245 3893 8248
rect 3927 8245 3939 8279
rect 3881 8239 3939 8245
rect 4893 8279 4951 8285
rect 4893 8245 4905 8279
rect 4939 8276 4951 8279
rect 5534 8276 5540 8288
rect 4939 8248 5540 8276
rect 4939 8245 4951 8248
rect 4893 8239 4951 8245
rect 5534 8236 5540 8248
rect 5592 8236 5598 8288
rect 1104 8186 5704 8208
rect 1104 8134 1753 8186
rect 1805 8134 1817 8186
rect 1869 8134 1881 8186
rect 1933 8134 1945 8186
rect 1997 8134 3294 8186
rect 3346 8134 3358 8186
rect 3410 8134 3422 8186
rect 3474 8134 3486 8186
rect 3538 8134 4836 8186
rect 4888 8134 4900 8186
rect 4952 8134 4964 8186
rect 5016 8134 5028 8186
rect 5080 8134 5704 8186
rect 1104 8112 5704 8134
rect 1578 8032 1584 8084
rect 1636 8072 1642 8084
rect 1765 8075 1823 8081
rect 1765 8072 1777 8075
rect 1636 8044 1777 8072
rect 1636 8032 1642 8044
rect 1765 8041 1777 8044
rect 1811 8041 1823 8075
rect 1765 8035 1823 8041
rect 4249 8007 4307 8013
rect 4249 7973 4261 8007
rect 4295 8004 4307 8007
rect 4430 8004 4436 8016
rect 4295 7976 4436 8004
rect 4295 7973 4307 7976
rect 4249 7967 4307 7973
rect 4430 7964 4436 7976
rect 4488 8004 4494 8016
rect 4801 8007 4859 8013
rect 4801 8004 4813 8007
rect 4488 7976 4813 8004
rect 4488 7964 4494 7976
rect 4801 7973 4813 7976
rect 4847 7973 4859 8007
rect 4801 7967 4859 7973
rect 2406 7828 2412 7880
rect 2464 7868 2470 7880
rect 2501 7871 2559 7877
rect 2501 7868 2513 7871
rect 2464 7840 2513 7868
rect 2464 7828 2470 7840
rect 2501 7837 2513 7840
rect 2547 7837 2559 7871
rect 2501 7831 2559 7837
rect 2777 7871 2835 7877
rect 2777 7837 2789 7871
rect 2823 7837 2835 7871
rect 2777 7831 2835 7837
rect 1486 7760 1492 7812
rect 1544 7800 1550 7812
rect 2792 7800 2820 7831
rect 3878 7828 3884 7880
rect 3936 7868 3942 7880
rect 3973 7871 4031 7877
rect 3973 7868 3985 7871
rect 3936 7840 3985 7868
rect 3936 7828 3942 7840
rect 3973 7837 3985 7840
rect 4019 7837 4031 7871
rect 3973 7831 4031 7837
rect 4062 7828 4068 7880
rect 4120 7868 4126 7880
rect 4341 7871 4399 7877
rect 4120 7840 4165 7868
rect 4120 7828 4126 7840
rect 4341 7837 4353 7871
rect 4387 7837 4399 7871
rect 4341 7831 4399 7837
rect 1544 7772 2820 7800
rect 1544 7760 1550 7772
rect 3602 7760 3608 7812
rect 3660 7800 3666 7812
rect 4356 7800 4384 7831
rect 4706 7828 4712 7880
rect 4764 7868 4770 7880
rect 4985 7871 5043 7877
rect 4985 7868 4997 7871
rect 4764 7840 4997 7868
rect 4764 7828 4770 7840
rect 4985 7837 4997 7840
rect 5031 7837 5043 7871
rect 4985 7831 5043 7837
rect 3660 7772 4384 7800
rect 3660 7760 3666 7772
rect 3786 7732 3792 7744
rect 3747 7704 3792 7732
rect 3786 7692 3792 7704
rect 3844 7692 3850 7744
rect 1104 7642 5704 7664
rect 1104 7590 2523 7642
rect 2575 7590 2587 7642
rect 2639 7590 2651 7642
rect 2703 7590 2715 7642
rect 2767 7590 4065 7642
rect 4117 7590 4129 7642
rect 4181 7590 4193 7642
rect 4245 7590 4257 7642
rect 4309 7590 5704 7642
rect 1104 7568 5704 7590
rect 2314 7488 2320 7540
rect 2372 7528 2378 7540
rect 2501 7531 2559 7537
rect 2501 7528 2513 7531
rect 2372 7500 2513 7528
rect 2372 7488 2378 7500
rect 2501 7497 2513 7500
rect 2547 7497 2559 7531
rect 2501 7491 2559 7497
rect 4157 7531 4215 7537
rect 4157 7497 4169 7531
rect 4203 7497 4215 7531
rect 4157 7491 4215 7497
rect 4172 7460 4200 7491
rect 3252 7432 4200 7460
rect 1765 7395 1823 7401
rect 1765 7361 1777 7395
rect 1811 7392 1823 7395
rect 2130 7392 2136 7404
rect 1811 7364 2136 7392
rect 1811 7361 1823 7364
rect 1765 7355 1823 7361
rect 2130 7352 2136 7364
rect 2188 7352 2194 7404
rect 3252 7401 3280 7432
rect 3237 7395 3295 7401
rect 3237 7361 3249 7395
rect 3283 7361 3295 7395
rect 3237 7355 3295 7361
rect 3421 7395 3479 7401
rect 3421 7361 3433 7395
rect 3467 7392 3479 7395
rect 3602 7392 3608 7404
rect 3467 7364 3608 7392
rect 3467 7361 3479 7364
rect 3421 7355 3479 7361
rect 3602 7352 3608 7364
rect 3660 7352 3666 7404
rect 3697 7395 3755 7401
rect 3697 7361 3709 7395
rect 3743 7361 3755 7395
rect 3697 7355 3755 7361
rect 1486 7324 1492 7336
rect 1447 7296 1492 7324
rect 1486 7284 1492 7296
rect 1544 7284 1550 7336
rect 3513 7259 3571 7265
rect 3513 7225 3525 7259
rect 3559 7256 3571 7259
rect 3602 7256 3608 7268
rect 3559 7228 3608 7256
rect 3559 7225 3571 7228
rect 3513 7219 3571 7225
rect 3602 7216 3608 7228
rect 3660 7216 3666 7268
rect 3712 7256 3740 7355
rect 3878 7352 3884 7404
rect 3936 7392 3942 7404
rect 4341 7395 4399 7401
rect 4341 7392 4353 7395
rect 3936 7364 4353 7392
rect 3936 7352 3942 7364
rect 4341 7361 4353 7364
rect 4387 7361 4399 7395
rect 4341 7355 4399 7361
rect 4801 7395 4859 7401
rect 4801 7361 4813 7395
rect 4847 7361 4859 7395
rect 4801 7355 4859 7361
rect 4522 7324 4528 7336
rect 4483 7296 4528 7324
rect 4522 7284 4528 7296
rect 4580 7284 4586 7336
rect 4706 7256 4712 7268
rect 3712 7228 4712 7256
rect 4706 7216 4712 7228
rect 4764 7256 4770 7268
rect 4816 7256 4844 7355
rect 4764 7228 4844 7256
rect 4764 7216 4770 7228
rect 2774 7148 2780 7200
rect 2832 7188 2838 7200
rect 2961 7191 3019 7197
rect 2961 7188 2973 7191
rect 2832 7160 2973 7188
rect 2832 7148 2838 7160
rect 2961 7157 2973 7160
rect 3007 7157 3019 7191
rect 2961 7151 3019 7157
rect 3329 7191 3387 7197
rect 3329 7157 3341 7191
rect 3375 7188 3387 7191
rect 3694 7188 3700 7200
rect 3375 7160 3700 7188
rect 3375 7157 3387 7160
rect 3329 7151 3387 7157
rect 3694 7148 3700 7160
rect 3752 7188 3758 7200
rect 4430 7188 4436 7200
rect 3752 7160 4436 7188
rect 3752 7148 3758 7160
rect 4430 7148 4436 7160
rect 4488 7148 4494 7200
rect 1104 7098 5704 7120
rect 1104 7046 1753 7098
rect 1805 7046 1817 7098
rect 1869 7046 1881 7098
rect 1933 7046 1945 7098
rect 1997 7046 3294 7098
rect 3346 7046 3358 7098
rect 3410 7046 3422 7098
rect 3474 7046 3486 7098
rect 3538 7046 4836 7098
rect 4888 7046 4900 7098
rect 4952 7046 4964 7098
rect 5016 7046 5028 7098
rect 5080 7046 5704 7098
rect 1104 7024 5704 7046
rect 2225 6987 2283 6993
rect 2225 6953 2237 6987
rect 2271 6984 2283 6987
rect 2406 6984 2412 6996
rect 2271 6956 2412 6984
rect 2271 6953 2283 6956
rect 2225 6947 2283 6953
rect 2406 6944 2412 6956
rect 2464 6944 2470 6996
rect 3602 6944 3608 6996
rect 3660 6984 3666 6996
rect 3973 6987 4031 6993
rect 3973 6984 3985 6987
rect 3660 6956 3985 6984
rect 3660 6944 3666 6956
rect 3973 6953 3985 6956
rect 4019 6984 4031 6987
rect 4430 6984 4436 6996
rect 4019 6956 4436 6984
rect 4019 6953 4031 6956
rect 3973 6947 4031 6953
rect 4430 6944 4436 6956
rect 4488 6944 4494 6996
rect 1578 6876 1584 6928
rect 1636 6916 1642 6928
rect 2961 6919 3019 6925
rect 2961 6916 2973 6919
rect 1636 6888 2973 6916
rect 1636 6876 1642 6888
rect 2961 6885 2973 6888
rect 3007 6885 3019 6919
rect 2961 6879 3019 6885
rect 3786 6876 3792 6928
rect 3844 6916 3850 6928
rect 3844 6888 4200 6916
rect 3844 6876 3850 6888
rect 2222 6848 2228 6860
rect 2183 6820 2228 6848
rect 2222 6808 2228 6820
rect 2280 6808 2286 6860
rect 2317 6851 2375 6857
rect 2317 6817 2329 6851
rect 2363 6848 2375 6851
rect 2774 6848 2780 6860
rect 2363 6820 2780 6848
rect 2363 6817 2375 6820
rect 2317 6811 2375 6817
rect 2774 6808 2780 6820
rect 2832 6808 2838 6860
rect 2869 6851 2927 6857
rect 2869 6817 2881 6851
rect 2915 6848 2927 6851
rect 3602 6848 3608 6860
rect 2915 6820 3608 6848
rect 2915 6817 2927 6820
rect 2869 6811 2927 6817
rect 3602 6808 3608 6820
rect 3660 6808 3666 6860
rect 1394 6780 1400 6792
rect 1355 6752 1400 6780
rect 1394 6740 1400 6752
rect 1452 6740 1458 6792
rect 2406 6780 2412 6792
rect 2367 6752 2412 6780
rect 2406 6740 2412 6752
rect 2464 6740 2470 6792
rect 3053 6783 3111 6789
rect 3053 6749 3065 6783
rect 3099 6749 3111 6783
rect 3053 6743 3111 6749
rect 2038 6712 2044 6724
rect 1999 6684 2044 6712
rect 2038 6672 2044 6684
rect 2096 6672 2102 6724
rect 2866 6672 2872 6724
rect 2924 6712 2930 6724
rect 3068 6712 3096 6743
rect 3142 6740 3148 6792
rect 3200 6780 3206 6792
rect 4172 6789 4200 6888
rect 4706 6848 4712 6860
rect 4264 6820 4712 6848
rect 4065 6783 4123 6789
rect 3200 6752 3245 6780
rect 3200 6740 3206 6752
rect 4065 6749 4077 6783
rect 4111 6749 4123 6783
rect 4065 6743 4123 6749
rect 4157 6783 4215 6789
rect 4157 6749 4169 6783
rect 4203 6749 4215 6783
rect 4157 6743 4215 6749
rect 2924 6684 3096 6712
rect 4080 6712 4108 6743
rect 4264 6712 4292 6820
rect 4706 6808 4712 6820
rect 4764 6808 4770 6860
rect 4614 6740 4620 6792
rect 4672 6780 4678 6792
rect 4893 6783 4951 6789
rect 4893 6780 4905 6783
rect 4672 6752 4905 6780
rect 4672 6740 4678 6752
rect 4893 6749 4905 6752
rect 4939 6749 4951 6783
rect 4893 6743 4951 6749
rect 4080 6684 4292 6712
rect 2924 6672 2930 6684
rect 1486 6604 1492 6656
rect 1544 6644 1550 6656
rect 1581 6647 1639 6653
rect 1581 6644 1593 6647
rect 1544 6616 1593 6644
rect 1544 6604 1550 6616
rect 1581 6613 1593 6616
rect 1627 6613 1639 6647
rect 1581 6607 1639 6613
rect 2958 6604 2964 6656
rect 3016 6644 3022 6656
rect 3789 6647 3847 6653
rect 3789 6644 3801 6647
rect 3016 6616 3801 6644
rect 3016 6604 3022 6616
rect 3789 6613 3801 6616
rect 3835 6613 3847 6647
rect 3789 6607 3847 6613
rect 4522 6604 4528 6656
rect 4580 6644 4586 6656
rect 4709 6647 4767 6653
rect 4709 6644 4721 6647
rect 4580 6616 4721 6644
rect 4580 6604 4586 6616
rect 4709 6613 4721 6616
rect 4755 6613 4767 6647
rect 4709 6607 4767 6613
rect 1104 6554 5704 6576
rect 1104 6502 2523 6554
rect 2575 6502 2587 6554
rect 2639 6502 2651 6554
rect 2703 6502 2715 6554
rect 2767 6502 4065 6554
rect 4117 6502 4129 6554
rect 4181 6502 4193 6554
rect 4245 6502 4257 6554
rect 4309 6502 5704 6554
rect 1104 6480 5704 6502
rect 2875 6443 2933 6449
rect 2875 6409 2887 6443
rect 2921 6440 2933 6443
rect 3142 6440 3148 6452
rect 2921 6412 3148 6440
rect 2921 6409 2933 6412
rect 2875 6403 2933 6409
rect 3142 6400 3148 6412
rect 3200 6400 3206 6452
rect 4706 6440 4712 6452
rect 4667 6412 4712 6440
rect 4706 6400 4712 6412
rect 4764 6400 4770 6452
rect 2019 6375 2077 6381
rect 2019 6341 2031 6375
rect 2065 6372 2077 6375
rect 2130 6372 2136 6384
rect 2065 6344 2136 6372
rect 2065 6341 2077 6344
rect 2019 6335 2077 6341
rect 2130 6332 2136 6344
rect 2188 6332 2194 6384
rect 2958 6372 2964 6384
rect 2240 6344 2964 6372
rect 2240 6245 2268 6344
rect 2958 6332 2964 6344
rect 3016 6332 3022 6384
rect 3694 6332 3700 6384
rect 3752 6372 3758 6384
rect 4065 6375 4123 6381
rect 4065 6372 4077 6375
rect 3752 6344 4077 6372
rect 3752 6332 3758 6344
rect 4065 6341 4077 6344
rect 4111 6341 4123 6375
rect 4724 6372 4752 6400
rect 4065 6335 4123 6341
rect 4264 6344 4752 6372
rect 2317 6307 2375 6313
rect 2317 6273 2329 6307
rect 2363 6304 2375 6307
rect 2406 6304 2412 6316
rect 2363 6276 2412 6304
rect 2363 6273 2375 6276
rect 2317 6267 2375 6273
rect 2406 6264 2412 6276
rect 2464 6304 2470 6316
rect 2777 6307 2835 6313
rect 2777 6304 2789 6307
rect 2464 6276 2789 6304
rect 2464 6264 2470 6276
rect 2777 6273 2789 6276
rect 2823 6304 2835 6307
rect 2823 6276 3004 6304
rect 2823 6273 2835 6276
rect 2777 6267 2835 6273
rect 2976 6248 3004 6276
rect 3050 6264 3056 6316
rect 3108 6304 3114 6316
rect 3789 6307 3847 6313
rect 3108 6276 3153 6304
rect 3108 6264 3114 6276
rect 3789 6273 3801 6307
rect 3835 6304 3847 6307
rect 3970 6304 3976 6316
rect 3835 6276 3976 6304
rect 3835 6273 3847 6276
rect 3789 6267 3847 6273
rect 3970 6264 3976 6276
rect 4028 6304 4034 6316
rect 4264 6304 4292 6344
rect 4028 6276 4292 6304
rect 4525 6307 4583 6313
rect 4028 6264 4034 6276
rect 4525 6273 4537 6307
rect 4571 6304 4583 6307
rect 4706 6304 4712 6316
rect 4571 6276 4712 6304
rect 4571 6273 4583 6276
rect 4525 6267 4583 6273
rect 4706 6264 4712 6276
rect 4764 6264 4770 6316
rect 2133 6239 2191 6245
rect 2133 6205 2145 6239
rect 2179 6205 2191 6239
rect 2133 6199 2191 6205
rect 2225 6239 2283 6245
rect 2225 6205 2237 6239
rect 2271 6205 2283 6239
rect 2225 6199 2283 6205
rect 1949 6171 2007 6177
rect 1949 6137 1961 6171
rect 1995 6168 2007 6171
rect 2038 6168 2044 6180
rect 1995 6140 2044 6168
rect 1995 6137 2007 6140
rect 1949 6131 2007 6137
rect 1964 6100 1992 6131
rect 2038 6128 2044 6140
rect 2096 6128 2102 6180
rect 2148 6168 2176 6199
rect 2958 6196 2964 6248
rect 3016 6196 3022 6248
rect 3878 6236 3884 6248
rect 3839 6208 3884 6236
rect 3878 6196 3884 6208
rect 3936 6196 3942 6248
rect 2406 6168 2412 6180
rect 2148 6140 2412 6168
rect 2406 6128 2412 6140
rect 2464 6128 2470 6180
rect 3605 6103 3663 6109
rect 3605 6100 3617 6103
rect 1964 6072 3617 6100
rect 3605 6069 3617 6072
rect 3651 6069 3663 6103
rect 3605 6063 3663 6069
rect 4065 6103 4123 6109
rect 4065 6069 4077 6103
rect 4111 6100 4123 6103
rect 4430 6100 4436 6112
rect 4111 6072 4436 6100
rect 4111 6069 4123 6072
rect 4065 6063 4123 6069
rect 4430 6060 4436 6072
rect 4488 6100 4494 6112
rect 4614 6100 4620 6112
rect 4488 6072 4620 6100
rect 4488 6060 4494 6072
rect 4614 6060 4620 6072
rect 4672 6060 4678 6112
rect 1104 6010 5704 6032
rect 1104 5958 1753 6010
rect 1805 5958 1817 6010
rect 1869 5958 1881 6010
rect 1933 5958 1945 6010
rect 1997 5958 3294 6010
rect 3346 5958 3358 6010
rect 3410 5958 3422 6010
rect 3474 5958 3486 6010
rect 3538 5958 4836 6010
rect 4888 5958 4900 6010
rect 4952 5958 4964 6010
rect 5016 5958 5028 6010
rect 5080 5958 5704 6010
rect 1104 5936 5704 5958
rect 1673 5899 1731 5905
rect 1673 5865 1685 5899
rect 1719 5896 1731 5899
rect 2866 5896 2872 5908
rect 1719 5868 2872 5896
rect 1719 5865 1731 5868
rect 1673 5859 1731 5865
rect 2866 5856 2872 5868
rect 2924 5856 2930 5908
rect 5813 5831 5871 5837
rect 5813 5797 5825 5831
rect 5859 5828 5871 5831
rect 6638 5828 6644 5840
rect 5859 5800 6644 5828
rect 5859 5797 5871 5800
rect 5813 5791 5871 5797
rect 6638 5788 6644 5800
rect 6696 5788 6702 5840
rect 1578 5720 1584 5772
rect 1636 5760 1642 5772
rect 2225 5763 2283 5769
rect 2225 5760 2237 5763
rect 1636 5732 2237 5760
rect 1636 5720 1642 5732
rect 2225 5729 2237 5732
rect 2271 5729 2283 5763
rect 3970 5760 3976 5772
rect 3931 5732 3976 5760
rect 2225 5723 2283 5729
rect 3970 5720 3976 5732
rect 4028 5720 4034 5772
rect 4341 5763 4399 5769
rect 4341 5729 4353 5763
rect 4387 5760 4399 5763
rect 4430 5760 4436 5772
rect 4387 5732 4436 5760
rect 4387 5729 4399 5732
rect 4341 5723 4399 5729
rect 4430 5720 4436 5732
rect 4488 5720 4494 5772
rect 1394 5692 1400 5704
rect 1355 5664 1400 5692
rect 1394 5652 1400 5664
rect 1452 5652 1458 5704
rect 1673 5695 1731 5701
rect 1673 5661 1685 5695
rect 1719 5692 1731 5695
rect 2038 5692 2044 5704
rect 1719 5664 2044 5692
rect 1719 5661 1731 5664
rect 1673 5655 1731 5661
rect 2038 5652 2044 5664
rect 2096 5652 2102 5704
rect 2501 5695 2559 5701
rect 2501 5661 2513 5695
rect 2547 5692 2559 5695
rect 3142 5692 3148 5704
rect 2547 5664 3148 5692
rect 2547 5661 2559 5664
rect 2501 5655 2559 5661
rect 3142 5652 3148 5664
rect 3200 5652 3206 5704
rect 4065 5695 4123 5701
rect 4065 5661 4077 5695
rect 4111 5692 4123 5695
rect 4614 5692 4620 5704
rect 4111 5664 4620 5692
rect 4111 5661 4123 5664
rect 4065 5655 4123 5661
rect 4614 5652 4620 5664
rect 4672 5652 4678 5704
rect 2314 5584 2320 5636
rect 2372 5624 2378 5636
rect 4433 5627 4491 5633
rect 2372 5596 3188 5624
rect 2372 5584 2378 5596
rect 3160 5568 3188 5596
rect 3252 5596 4292 5624
rect 1489 5559 1547 5565
rect 1489 5525 1501 5559
rect 1535 5556 1547 5559
rect 2406 5556 2412 5568
rect 1535 5528 2412 5556
rect 1535 5525 1547 5528
rect 1489 5519 1547 5525
rect 2406 5516 2412 5528
rect 2464 5516 2470 5568
rect 3142 5516 3148 5568
rect 3200 5516 3206 5568
rect 3252 5565 3280 5596
rect 3237 5559 3295 5565
rect 3237 5525 3249 5559
rect 3283 5525 3295 5559
rect 3786 5556 3792 5568
rect 3747 5528 3792 5556
rect 3237 5519 3295 5525
rect 3786 5516 3792 5528
rect 3844 5516 3850 5568
rect 4264 5556 4292 5596
rect 4433 5593 4445 5627
rect 4479 5624 4491 5627
rect 4706 5624 4712 5636
rect 4479 5596 4712 5624
rect 4479 5593 4491 5596
rect 4433 5587 4491 5593
rect 4706 5584 4712 5596
rect 4764 5584 4770 5636
rect 4798 5556 4804 5568
rect 4264 5528 4804 5556
rect 4798 5516 4804 5528
rect 4856 5516 4862 5568
rect 1104 5466 5704 5488
rect 1104 5414 2523 5466
rect 2575 5414 2587 5466
rect 2639 5414 2651 5466
rect 2703 5414 2715 5466
rect 2767 5414 4065 5466
rect 4117 5414 4129 5466
rect 4181 5414 4193 5466
rect 4245 5414 4257 5466
rect 4309 5414 5704 5466
rect 1104 5392 5704 5414
rect 2406 5352 2412 5364
rect 2367 5324 2412 5352
rect 2406 5312 2412 5324
rect 2464 5312 2470 5364
rect 3050 5312 3056 5364
rect 3108 5352 3114 5364
rect 3605 5355 3663 5361
rect 3605 5352 3617 5355
rect 3108 5324 3617 5352
rect 3108 5312 3114 5324
rect 3605 5321 3617 5324
rect 3651 5321 3663 5355
rect 3605 5315 3663 5321
rect 1397 5287 1455 5293
rect 1397 5253 1409 5287
rect 1443 5284 1455 5287
rect 2590 5284 2596 5296
rect 1443 5256 2596 5284
rect 1443 5253 1455 5256
rect 1397 5247 1455 5253
rect 2590 5244 2596 5256
rect 2648 5244 2654 5296
rect 4798 5284 4804 5296
rect 4759 5256 4804 5284
rect 4798 5244 4804 5256
rect 4856 5244 4862 5296
rect 1486 5176 1492 5228
rect 1544 5216 1550 5228
rect 1581 5219 1639 5225
rect 1581 5216 1593 5219
rect 1544 5188 1593 5216
rect 1544 5176 1550 5188
rect 1581 5185 1593 5188
rect 1627 5185 1639 5219
rect 1581 5179 1639 5185
rect 1765 5219 1823 5225
rect 1765 5185 1777 5219
rect 1811 5216 1823 5219
rect 2130 5216 2136 5228
rect 1811 5188 2136 5216
rect 1811 5185 1823 5188
rect 1765 5179 1823 5185
rect 1596 5148 1624 5179
rect 2130 5176 2136 5188
rect 2188 5176 2194 5228
rect 2774 5216 2780 5228
rect 2735 5188 2780 5216
rect 2774 5176 2780 5188
rect 2832 5176 2838 5228
rect 3786 5176 3792 5228
rect 3844 5216 3850 5228
rect 3973 5219 4031 5225
rect 3973 5216 3985 5219
rect 3844 5188 3985 5216
rect 3844 5176 3850 5188
rect 3973 5185 3985 5188
rect 4019 5185 4031 5219
rect 3973 5179 4031 5185
rect 3050 5148 3056 5160
rect 1596 5120 3056 5148
rect 3050 5108 3056 5120
rect 3108 5108 3114 5160
rect 3878 5148 3884 5160
rect 3839 5120 3884 5148
rect 3878 5108 3884 5120
rect 3936 5108 3942 5160
rect 4985 5083 5043 5089
rect 4985 5049 4997 5083
rect 5031 5080 5043 5083
rect 5350 5080 5356 5092
rect 5031 5052 5356 5080
rect 5031 5049 5043 5052
rect 4985 5043 5043 5049
rect 5350 5040 5356 5052
rect 5408 5040 5414 5092
rect 3694 4972 3700 5024
rect 3752 5012 3758 5024
rect 3789 5015 3847 5021
rect 3789 5012 3801 5015
rect 3752 4984 3801 5012
rect 3752 4972 3758 4984
rect 3789 4981 3801 4984
rect 3835 4981 3847 5015
rect 3789 4975 3847 4981
rect 1104 4922 5704 4944
rect 1104 4870 1753 4922
rect 1805 4870 1817 4922
rect 1869 4870 1881 4922
rect 1933 4870 1945 4922
rect 1997 4870 3294 4922
rect 3346 4870 3358 4922
rect 3410 4870 3422 4922
rect 3474 4870 3486 4922
rect 3538 4870 4836 4922
rect 4888 4870 4900 4922
rect 4952 4870 4964 4922
rect 5016 4870 5028 4922
rect 5080 4870 5704 4922
rect 1104 4848 5704 4870
rect 1394 4808 1400 4820
rect 1355 4780 1400 4808
rect 1394 4768 1400 4780
rect 1452 4768 1458 4820
rect 2593 4811 2651 4817
rect 2593 4808 2605 4811
rect 1780 4780 2605 4808
rect 1780 4616 1808 4780
rect 2593 4777 2605 4780
rect 2639 4777 2651 4811
rect 2593 4771 2651 4777
rect 2774 4768 2780 4820
rect 2832 4808 2838 4820
rect 3789 4811 3847 4817
rect 3789 4808 3801 4811
rect 2832 4780 3801 4808
rect 2832 4768 2838 4780
rect 3789 4777 3801 4780
rect 3835 4777 3847 4811
rect 3789 4771 3847 4777
rect 2958 4740 2964 4752
rect 2919 4712 2964 4740
rect 2958 4700 2964 4712
rect 3016 4700 3022 4752
rect 1857 4675 1915 4681
rect 1857 4641 1869 4675
rect 1903 4672 1915 4675
rect 2685 4675 2743 4681
rect 2685 4672 2697 4675
rect 1903 4644 2697 4672
rect 1903 4641 1915 4644
rect 1857 4635 1915 4641
rect 2685 4641 2697 4644
rect 2731 4672 2743 4675
rect 2866 4672 2872 4684
rect 2731 4644 2872 4672
rect 2731 4641 2743 4644
rect 2685 4635 2743 4641
rect 2866 4632 2872 4644
rect 2924 4632 2930 4684
rect 4433 4675 4491 4681
rect 4433 4641 4445 4675
rect 4479 4672 4491 4675
rect 4522 4672 4528 4684
rect 4479 4644 4528 4672
rect 4479 4641 4491 4644
rect 4433 4635 4491 4641
rect 4522 4632 4528 4644
rect 4580 4632 4586 4684
rect 1578 4564 1584 4616
rect 1636 4604 1642 4616
rect 1673 4607 1731 4613
rect 1673 4604 1685 4607
rect 1636 4576 1685 4604
rect 1636 4564 1642 4576
rect 1673 4573 1685 4576
rect 1719 4573 1731 4607
rect 1673 4567 1731 4573
rect 1762 4564 1768 4616
rect 1820 4604 1826 4616
rect 2130 4604 2136 4616
rect 1820 4576 1865 4604
rect 2091 4576 2136 4604
rect 1820 4564 1826 4576
rect 2130 4564 2136 4576
rect 2188 4564 2194 4616
rect 2590 4604 2596 4616
rect 2551 4576 2596 4604
rect 2590 4564 2596 4576
rect 2648 4564 2654 4616
rect 2884 4604 2912 4632
rect 3914 4607 3972 4613
rect 3914 4604 3926 4607
rect 2884 4576 3926 4604
rect 3914 4573 3926 4576
rect 3960 4573 3972 4607
rect 3914 4567 3972 4573
rect 4341 4607 4399 4613
rect 4341 4573 4353 4607
rect 4387 4573 4399 4607
rect 4341 4567 4399 4573
rect 2041 4471 2099 4477
rect 2041 4437 2053 4471
rect 2087 4468 2099 4471
rect 2958 4468 2964 4480
rect 2087 4440 2964 4468
rect 2087 4437 2099 4440
rect 2041 4431 2099 4437
rect 2958 4428 2964 4440
rect 3016 4428 3022 4480
rect 3878 4428 3884 4480
rect 3936 4468 3942 4480
rect 3973 4471 4031 4477
rect 3973 4468 3985 4471
rect 3936 4440 3985 4468
rect 3936 4428 3942 4440
rect 3973 4437 3985 4440
rect 4019 4468 4031 4471
rect 4356 4468 4384 4567
rect 4019 4440 4384 4468
rect 4019 4437 4031 4440
rect 3973 4431 4031 4437
rect 1104 4378 5704 4400
rect 1104 4326 2523 4378
rect 2575 4326 2587 4378
rect 2639 4326 2651 4378
rect 2703 4326 2715 4378
rect 2767 4326 4065 4378
rect 4117 4326 4129 4378
rect 4181 4326 4193 4378
rect 4245 4326 4257 4378
rect 4309 4326 5704 4378
rect 1104 4304 5704 4326
rect 2866 4224 2872 4276
rect 2924 4264 2930 4276
rect 3513 4267 3571 4273
rect 3513 4264 3525 4267
rect 2924 4236 3525 4264
rect 2924 4224 2930 4236
rect 3513 4233 3525 4236
rect 3559 4233 3571 4267
rect 3513 4227 3571 4233
rect 4433 4267 4491 4273
rect 4433 4233 4445 4267
rect 4479 4264 4491 4267
rect 4614 4264 4620 4276
rect 4479 4236 4620 4264
rect 4479 4233 4491 4236
rect 4433 4227 4491 4233
rect 4614 4224 4620 4236
rect 4672 4224 4678 4276
rect 2130 4128 2136 4140
rect 2091 4100 2136 4128
rect 2130 4088 2136 4100
rect 2188 4088 2194 4140
rect 2593 4131 2651 4137
rect 2593 4097 2605 4131
rect 2639 4128 2651 4131
rect 2866 4128 2872 4140
rect 2639 4100 2872 4128
rect 2639 4097 2651 4100
rect 2593 4091 2651 4097
rect 2866 4088 2872 4100
rect 2924 4088 2930 4140
rect 3697 4131 3755 4137
rect 3697 4097 3709 4131
rect 3743 4097 3755 4131
rect 3697 4091 3755 4097
rect 4249 4131 4307 4137
rect 4249 4097 4261 4131
rect 4295 4128 4307 4131
rect 4430 4128 4436 4140
rect 4295 4100 4436 4128
rect 4295 4097 4307 4100
rect 4249 4091 4307 4097
rect 1857 4063 1915 4069
rect 1857 4029 1869 4063
rect 1903 4060 1915 4063
rect 2222 4060 2228 4072
rect 1903 4032 2228 4060
rect 1903 4029 1915 4032
rect 1857 4023 1915 4029
rect 2222 4020 2228 4032
rect 2280 4020 2286 4072
rect 3712 4060 3740 4091
rect 4430 4088 4436 4100
rect 4488 4088 4494 4140
rect 4522 4060 4528 4072
rect 3712 4032 4528 4060
rect 4522 4020 4528 4032
rect 4580 4020 4586 4072
rect 1762 3952 1768 4004
rect 1820 3992 1826 4004
rect 2409 3995 2467 4001
rect 2409 3992 2421 3995
rect 1820 3964 2421 3992
rect 1820 3952 1826 3964
rect 2409 3961 2421 3964
rect 2455 3992 2467 3995
rect 2498 3992 2504 4004
rect 2455 3964 2504 3992
rect 2455 3961 2467 3964
rect 2409 3955 2467 3961
rect 2498 3952 2504 3964
rect 2556 3952 2562 4004
rect 2038 3884 2044 3936
rect 2096 3924 2102 3936
rect 2225 3927 2283 3933
rect 2225 3924 2237 3927
rect 2096 3896 2237 3924
rect 2096 3884 2102 3896
rect 2225 3893 2237 3896
rect 2271 3893 2283 3927
rect 2225 3887 2283 3893
rect 2314 3884 2320 3936
rect 2372 3924 2378 3936
rect 2372 3896 2417 3924
rect 2372 3884 2378 3896
rect 1104 3834 5704 3856
rect 1104 3782 1753 3834
rect 1805 3782 1817 3834
rect 1869 3782 1881 3834
rect 1933 3782 1945 3834
rect 1997 3782 3294 3834
rect 3346 3782 3358 3834
rect 3410 3782 3422 3834
rect 3474 3782 3486 3834
rect 3538 3782 4836 3834
rect 4888 3782 4900 3834
rect 4952 3782 4964 3834
rect 5016 3782 5028 3834
rect 5080 3782 5704 3834
rect 1104 3760 5704 3782
rect 1578 3720 1584 3732
rect 1539 3692 1584 3720
rect 1578 3680 1584 3692
rect 1636 3680 1642 3732
rect 2130 3720 2136 3732
rect 2091 3692 2136 3720
rect 2130 3680 2136 3692
rect 2188 3680 2194 3732
rect 2222 3680 2228 3732
rect 2280 3720 2286 3732
rect 2317 3723 2375 3729
rect 2317 3720 2329 3723
rect 2280 3692 2329 3720
rect 2280 3680 2286 3692
rect 2317 3689 2329 3692
rect 2363 3720 2375 3723
rect 2498 3720 2504 3732
rect 2363 3692 2504 3720
rect 2363 3689 2375 3692
rect 2317 3683 2375 3689
rect 2498 3680 2504 3692
rect 2556 3680 2562 3732
rect 3878 3720 3884 3732
rect 3839 3692 3884 3720
rect 3878 3680 3884 3692
rect 3936 3680 3942 3732
rect 4801 3723 4859 3729
rect 4801 3689 4813 3723
rect 4847 3720 4859 3723
rect 5905 3723 5963 3729
rect 5905 3720 5917 3723
rect 4847 3692 5917 3720
rect 4847 3689 4859 3692
rect 4801 3683 4859 3689
rect 5905 3689 5917 3692
rect 5951 3689 5963 3723
rect 5905 3683 5963 3689
rect 2406 3584 2412 3596
rect 1504 3556 2412 3584
rect 1504 3525 1532 3556
rect 2406 3544 2412 3556
rect 2464 3544 2470 3596
rect 2516 3584 2544 3680
rect 2516 3556 3832 3584
rect 1489 3519 1547 3525
rect 1489 3485 1501 3519
rect 1535 3485 1547 3519
rect 1489 3479 1547 3485
rect 2685 3519 2743 3525
rect 2685 3485 2697 3519
rect 2731 3516 2743 3519
rect 2866 3516 2872 3528
rect 2731 3488 2872 3516
rect 2731 3485 2743 3488
rect 2685 3479 2743 3485
rect 2866 3476 2872 3488
rect 2924 3476 2930 3528
rect 3804 3525 3832 3556
rect 3789 3519 3847 3525
rect 3789 3485 3801 3519
rect 3835 3485 3847 3519
rect 3789 3479 3847 3485
rect 4985 3519 5043 3525
rect 4985 3485 4997 3519
rect 5031 3516 5043 3519
rect 5813 3519 5871 3525
rect 5813 3516 5825 3519
rect 5031 3488 5825 3516
rect 5031 3485 5043 3488
rect 4985 3479 5043 3485
rect 5813 3485 5825 3488
rect 5859 3485 5871 3519
rect 5813 3479 5871 3485
rect 1104 3290 5704 3312
rect 1104 3238 2523 3290
rect 2575 3238 2587 3290
rect 2639 3238 2651 3290
rect 2703 3238 2715 3290
rect 2767 3238 4065 3290
rect 4117 3238 4129 3290
rect 4181 3238 4193 3290
rect 4245 3238 4257 3290
rect 4309 3238 5704 3290
rect 1104 3216 5704 3238
rect 1581 3179 1639 3185
rect 1581 3145 1593 3179
rect 1627 3176 1639 3179
rect 2038 3176 2044 3188
rect 1627 3148 2044 3176
rect 1627 3145 1639 3148
rect 1581 3139 1639 3145
rect 2038 3136 2044 3148
rect 2096 3136 2102 3188
rect 2314 3136 2320 3188
rect 2372 3176 2378 3188
rect 2869 3179 2927 3185
rect 2869 3176 2881 3179
rect 2372 3148 2881 3176
rect 2372 3136 2378 3148
rect 2869 3145 2881 3148
rect 2915 3145 2927 3179
rect 2869 3139 2927 3145
rect 3605 3179 3663 3185
rect 3605 3145 3617 3179
rect 3651 3145 3663 3179
rect 3605 3139 3663 3145
rect 3620 3108 3648 3139
rect 3786 3136 3792 3188
rect 3844 3176 3850 3188
rect 4341 3179 4399 3185
rect 4341 3176 4353 3179
rect 3844 3148 4353 3176
rect 3844 3136 3850 3148
rect 4341 3145 4353 3148
rect 4387 3145 4399 3179
rect 4341 3139 4399 3145
rect 4706 3108 4712 3120
rect 3620 3080 4712 3108
rect 4706 3068 4712 3080
rect 4764 3068 4770 3120
rect 1394 3040 1400 3052
rect 1355 3012 1400 3040
rect 1394 3000 1400 3012
rect 1452 3000 1458 3052
rect 2038 3000 2044 3052
rect 2096 3040 2102 3052
rect 2133 3043 2191 3049
rect 2133 3040 2145 3043
rect 2096 3012 2145 3040
rect 2096 3000 2102 3012
rect 2133 3009 2145 3012
rect 2179 3009 2191 3043
rect 2133 3003 2191 3009
rect 2317 3043 2375 3049
rect 2317 3009 2329 3043
rect 2363 3009 2375 3043
rect 2317 3003 2375 3009
rect 2777 3043 2835 3049
rect 2777 3009 2789 3043
rect 2823 3040 2835 3043
rect 2958 3040 2964 3052
rect 2823 3012 2964 3040
rect 2823 3009 2835 3012
rect 2777 3003 2835 3009
rect 2332 2972 2360 3003
rect 2958 3000 2964 3012
rect 3016 3000 3022 3052
rect 3142 3000 3148 3052
rect 3200 3040 3206 3052
rect 3421 3043 3479 3049
rect 3421 3040 3433 3043
rect 3200 3012 3433 3040
rect 3200 3000 3206 3012
rect 3421 3009 3433 3012
rect 3467 3009 3479 3043
rect 3421 3003 3479 3009
rect 3878 3000 3884 3052
rect 3936 3040 3942 3052
rect 4157 3043 4215 3049
rect 4157 3040 4169 3043
rect 3936 3012 4169 3040
rect 3936 3000 3942 3012
rect 4157 3009 4169 3012
rect 4203 3009 4215 3043
rect 4157 3003 4215 3009
rect 4801 3043 4859 3049
rect 4801 3009 4813 3043
rect 4847 3040 4859 3043
rect 5997 3043 6055 3049
rect 5997 3040 6009 3043
rect 4847 3012 6009 3040
rect 4847 3009 4859 3012
rect 4801 3003 4859 3009
rect 5997 3009 6009 3012
rect 6043 3009 6055 3043
rect 5997 3003 6055 3009
rect 2866 2972 2872 2984
rect 2332 2944 2872 2972
rect 2866 2932 2872 2944
rect 2924 2932 2930 2984
rect 2225 2907 2283 2913
rect 2225 2873 2237 2907
rect 2271 2904 2283 2907
rect 4816 2904 4844 3003
rect 2271 2876 4844 2904
rect 2271 2873 2283 2876
rect 2225 2867 2283 2873
rect 4706 2796 4712 2848
rect 4764 2836 4770 2848
rect 4893 2839 4951 2845
rect 4893 2836 4905 2839
rect 4764 2808 4905 2836
rect 4764 2796 4770 2808
rect 4893 2805 4905 2808
rect 4939 2805 4951 2839
rect 4893 2799 4951 2805
rect 1104 2746 5704 2768
rect 1104 2694 1753 2746
rect 1805 2694 1817 2746
rect 1869 2694 1881 2746
rect 1933 2694 1945 2746
rect 1997 2694 3294 2746
rect 3346 2694 3358 2746
rect 3410 2694 3422 2746
rect 3474 2694 3486 2746
rect 3538 2694 4836 2746
rect 4888 2694 4900 2746
rect 4952 2694 4964 2746
rect 5016 2694 5028 2746
rect 5080 2694 5704 2746
rect 1104 2672 5704 2694
rect 2866 2632 2872 2644
rect 2779 2604 2872 2632
rect 2866 2592 2872 2604
rect 2924 2632 2930 2644
rect 3602 2632 3608 2644
rect 2924 2604 3608 2632
rect 2924 2592 2930 2604
rect 3602 2592 3608 2604
rect 3660 2592 3666 2644
rect 4249 2635 4307 2641
rect 4249 2601 4261 2635
rect 4295 2632 4307 2635
rect 4430 2632 4436 2644
rect 4295 2604 4436 2632
rect 4295 2601 4307 2604
rect 4249 2595 4307 2601
rect 4430 2592 4436 2604
rect 4488 2592 4494 2644
rect 1673 2499 1731 2505
rect 1673 2465 1685 2499
rect 1719 2496 1731 2499
rect 2222 2496 2228 2508
rect 1719 2468 2228 2496
rect 1719 2465 1731 2468
rect 1673 2459 1731 2465
rect 2222 2456 2228 2468
rect 2280 2456 2286 2508
rect 14 2388 20 2440
rect 72 2428 78 2440
rect 1397 2431 1455 2437
rect 1397 2428 1409 2431
rect 72 2400 1409 2428
rect 72 2388 78 2400
rect 1397 2397 1409 2400
rect 1443 2397 1455 2431
rect 1397 2391 1455 2397
rect 2038 2388 2044 2440
rect 2096 2428 2102 2440
rect 2685 2431 2743 2437
rect 2685 2428 2697 2431
rect 2096 2400 2697 2428
rect 2096 2388 2102 2400
rect 2685 2397 2697 2400
rect 2731 2397 2743 2431
rect 4062 2428 4068 2440
rect 4023 2400 4068 2428
rect 2685 2391 2743 2397
rect 4062 2388 4068 2400
rect 4120 2388 4126 2440
rect 4706 2388 4712 2440
rect 4764 2428 4770 2440
rect 4801 2431 4859 2437
rect 4801 2428 4813 2431
rect 4764 2400 4813 2428
rect 4764 2388 4770 2400
rect 4801 2397 4813 2400
rect 4847 2397 4859 2431
rect 4801 2391 4859 2397
rect 4985 2363 5043 2369
rect 4985 2329 4997 2363
rect 5031 2360 5043 2363
rect 6086 2360 6092 2372
rect 5031 2332 6092 2360
rect 5031 2329 5043 2332
rect 4985 2323 5043 2329
rect 6086 2320 6092 2332
rect 6144 2320 6150 2372
rect 1104 2202 5704 2224
rect 1104 2150 2523 2202
rect 2575 2150 2587 2202
rect 2639 2150 2651 2202
rect 2703 2150 2715 2202
rect 2767 2150 4065 2202
rect 4117 2150 4129 2202
rect 4181 2150 4193 2202
rect 4245 2150 4257 2202
rect 4309 2150 5704 2202
rect 1104 2128 5704 2150
<< via1 >>
rect 2523 8678 2575 8730
rect 2587 8678 2639 8730
rect 2651 8678 2703 8730
rect 2715 8678 2767 8730
rect 4065 8678 4117 8730
rect 4129 8678 4181 8730
rect 4193 8678 4245 8730
rect 4257 8678 4309 8730
rect 1492 8619 1544 8628
rect 1492 8585 1501 8619
rect 1501 8585 1535 8619
rect 1535 8585 1544 8619
rect 1492 8576 1544 8585
rect 572 8508 624 8560
rect 1584 8483 1636 8492
rect 1584 8449 1593 8483
rect 1593 8449 1627 8483
rect 1627 8449 1636 8483
rect 1584 8440 1636 8449
rect 2320 8483 2372 8492
rect 2320 8449 2329 8483
rect 2329 8449 2363 8483
rect 2363 8449 2372 8483
rect 2320 8440 2372 8449
rect 3884 8440 3936 8492
rect 4712 8372 4764 8424
rect 4068 8304 4120 8356
rect 3608 8236 3660 8288
rect 5540 8236 5592 8288
rect 1753 8134 1805 8186
rect 1817 8134 1869 8186
rect 1881 8134 1933 8186
rect 1945 8134 1997 8186
rect 3294 8134 3346 8186
rect 3358 8134 3410 8186
rect 3422 8134 3474 8186
rect 3486 8134 3538 8186
rect 4836 8134 4888 8186
rect 4900 8134 4952 8186
rect 4964 8134 5016 8186
rect 5028 8134 5080 8186
rect 1584 8032 1636 8084
rect 4436 7964 4488 8016
rect 2412 7828 2464 7880
rect 1492 7760 1544 7812
rect 3884 7828 3936 7880
rect 4068 7871 4120 7880
rect 4068 7837 4077 7871
rect 4077 7837 4111 7871
rect 4111 7837 4120 7871
rect 4068 7828 4120 7837
rect 3608 7760 3660 7812
rect 4712 7828 4764 7880
rect 3792 7735 3844 7744
rect 3792 7701 3801 7735
rect 3801 7701 3835 7735
rect 3835 7701 3844 7735
rect 3792 7692 3844 7701
rect 2523 7590 2575 7642
rect 2587 7590 2639 7642
rect 2651 7590 2703 7642
rect 2715 7590 2767 7642
rect 4065 7590 4117 7642
rect 4129 7590 4181 7642
rect 4193 7590 4245 7642
rect 4257 7590 4309 7642
rect 2320 7488 2372 7540
rect 2136 7352 2188 7404
rect 3608 7352 3660 7404
rect 1492 7327 1544 7336
rect 1492 7293 1501 7327
rect 1501 7293 1535 7327
rect 1535 7293 1544 7327
rect 1492 7284 1544 7293
rect 3608 7216 3660 7268
rect 3884 7352 3936 7404
rect 4528 7327 4580 7336
rect 4528 7293 4537 7327
rect 4537 7293 4571 7327
rect 4571 7293 4580 7327
rect 4528 7284 4580 7293
rect 4712 7216 4764 7268
rect 2780 7148 2832 7200
rect 3700 7148 3752 7200
rect 4436 7191 4488 7200
rect 4436 7157 4445 7191
rect 4445 7157 4479 7191
rect 4479 7157 4488 7191
rect 4436 7148 4488 7157
rect 1753 7046 1805 7098
rect 1817 7046 1869 7098
rect 1881 7046 1933 7098
rect 1945 7046 1997 7098
rect 3294 7046 3346 7098
rect 3358 7046 3410 7098
rect 3422 7046 3474 7098
rect 3486 7046 3538 7098
rect 4836 7046 4888 7098
rect 4900 7046 4952 7098
rect 4964 7046 5016 7098
rect 5028 7046 5080 7098
rect 2412 6944 2464 6996
rect 3608 6944 3660 6996
rect 4436 6944 4488 6996
rect 1584 6876 1636 6928
rect 3792 6876 3844 6928
rect 2228 6851 2280 6860
rect 2228 6817 2237 6851
rect 2237 6817 2271 6851
rect 2271 6817 2280 6851
rect 2228 6808 2280 6817
rect 2780 6808 2832 6860
rect 3608 6808 3660 6860
rect 1400 6783 1452 6792
rect 1400 6749 1409 6783
rect 1409 6749 1443 6783
rect 1443 6749 1452 6783
rect 1400 6740 1452 6749
rect 2412 6783 2464 6792
rect 2412 6749 2421 6783
rect 2421 6749 2455 6783
rect 2455 6749 2464 6783
rect 2412 6740 2464 6749
rect 2044 6715 2096 6724
rect 2044 6681 2053 6715
rect 2053 6681 2087 6715
rect 2087 6681 2096 6715
rect 2044 6672 2096 6681
rect 2872 6672 2924 6724
rect 3148 6783 3200 6792
rect 3148 6749 3157 6783
rect 3157 6749 3191 6783
rect 3191 6749 3200 6783
rect 3148 6740 3200 6749
rect 4712 6808 4764 6860
rect 4620 6740 4672 6792
rect 1492 6604 1544 6656
rect 2964 6604 3016 6656
rect 4528 6604 4580 6656
rect 2523 6502 2575 6554
rect 2587 6502 2639 6554
rect 2651 6502 2703 6554
rect 2715 6502 2767 6554
rect 4065 6502 4117 6554
rect 4129 6502 4181 6554
rect 4193 6502 4245 6554
rect 4257 6502 4309 6554
rect 3148 6400 3200 6452
rect 4712 6443 4764 6452
rect 4712 6409 4721 6443
rect 4721 6409 4755 6443
rect 4755 6409 4764 6443
rect 4712 6400 4764 6409
rect 2136 6332 2188 6384
rect 2964 6375 3016 6384
rect 2964 6341 2973 6375
rect 2973 6341 3007 6375
rect 3007 6341 3016 6375
rect 2964 6332 3016 6341
rect 3700 6332 3752 6384
rect 2412 6264 2464 6316
rect 3056 6307 3108 6316
rect 3056 6273 3065 6307
rect 3065 6273 3099 6307
rect 3099 6273 3108 6307
rect 3056 6264 3108 6273
rect 3976 6264 4028 6316
rect 4712 6264 4764 6316
rect 2044 6128 2096 6180
rect 2964 6196 3016 6248
rect 3884 6239 3936 6248
rect 3884 6205 3893 6239
rect 3893 6205 3927 6239
rect 3927 6205 3936 6239
rect 3884 6196 3936 6205
rect 2412 6128 2464 6180
rect 4436 6060 4488 6112
rect 4620 6060 4672 6112
rect 1753 5958 1805 6010
rect 1817 5958 1869 6010
rect 1881 5958 1933 6010
rect 1945 5958 1997 6010
rect 3294 5958 3346 6010
rect 3358 5958 3410 6010
rect 3422 5958 3474 6010
rect 3486 5958 3538 6010
rect 4836 5958 4888 6010
rect 4900 5958 4952 6010
rect 4964 5958 5016 6010
rect 5028 5958 5080 6010
rect 2872 5856 2924 5908
rect 6644 5788 6696 5840
rect 1584 5720 1636 5772
rect 3976 5763 4028 5772
rect 3976 5729 3985 5763
rect 3985 5729 4019 5763
rect 4019 5729 4028 5763
rect 3976 5720 4028 5729
rect 4436 5720 4488 5772
rect 1400 5695 1452 5704
rect 1400 5661 1409 5695
rect 1409 5661 1443 5695
rect 1443 5661 1452 5695
rect 1400 5652 1452 5661
rect 2044 5652 2096 5704
rect 3148 5652 3200 5704
rect 4620 5652 4672 5704
rect 2320 5584 2372 5636
rect 2412 5516 2464 5568
rect 3148 5516 3200 5568
rect 3792 5559 3844 5568
rect 3792 5525 3801 5559
rect 3801 5525 3835 5559
rect 3835 5525 3844 5559
rect 3792 5516 3844 5525
rect 4712 5584 4764 5636
rect 4804 5516 4856 5568
rect 2523 5414 2575 5466
rect 2587 5414 2639 5466
rect 2651 5414 2703 5466
rect 2715 5414 2767 5466
rect 4065 5414 4117 5466
rect 4129 5414 4181 5466
rect 4193 5414 4245 5466
rect 4257 5414 4309 5466
rect 2412 5355 2464 5364
rect 2412 5321 2421 5355
rect 2421 5321 2455 5355
rect 2455 5321 2464 5355
rect 2412 5312 2464 5321
rect 3056 5312 3108 5364
rect 2596 5287 2648 5296
rect 2596 5253 2605 5287
rect 2605 5253 2639 5287
rect 2639 5253 2648 5287
rect 2596 5244 2648 5253
rect 4804 5287 4856 5296
rect 4804 5253 4813 5287
rect 4813 5253 4847 5287
rect 4847 5253 4856 5287
rect 4804 5244 4856 5253
rect 1492 5176 1544 5228
rect 2136 5176 2188 5228
rect 2780 5219 2832 5228
rect 2780 5185 2789 5219
rect 2789 5185 2823 5219
rect 2823 5185 2832 5219
rect 2780 5176 2832 5185
rect 3792 5176 3844 5228
rect 3056 5108 3108 5160
rect 3884 5151 3936 5160
rect 3884 5117 3893 5151
rect 3893 5117 3927 5151
rect 3927 5117 3936 5151
rect 3884 5108 3936 5117
rect 5356 5040 5408 5092
rect 3700 4972 3752 5024
rect 1753 4870 1805 4922
rect 1817 4870 1869 4922
rect 1881 4870 1933 4922
rect 1945 4870 1997 4922
rect 3294 4870 3346 4922
rect 3358 4870 3410 4922
rect 3422 4870 3474 4922
rect 3486 4870 3538 4922
rect 4836 4870 4888 4922
rect 4900 4870 4952 4922
rect 4964 4870 5016 4922
rect 5028 4870 5080 4922
rect 1400 4811 1452 4820
rect 1400 4777 1409 4811
rect 1409 4777 1443 4811
rect 1443 4777 1452 4811
rect 1400 4768 1452 4777
rect 2780 4768 2832 4820
rect 2964 4743 3016 4752
rect 2964 4709 2973 4743
rect 2973 4709 3007 4743
rect 3007 4709 3016 4743
rect 2964 4700 3016 4709
rect 2872 4632 2924 4684
rect 4528 4632 4580 4684
rect 1584 4564 1636 4616
rect 1768 4607 1820 4616
rect 1768 4573 1777 4607
rect 1777 4573 1811 4607
rect 1811 4573 1820 4607
rect 2136 4607 2188 4616
rect 1768 4564 1820 4573
rect 2136 4573 2145 4607
rect 2145 4573 2179 4607
rect 2179 4573 2188 4607
rect 2136 4564 2188 4573
rect 2596 4607 2648 4616
rect 2596 4573 2605 4607
rect 2605 4573 2639 4607
rect 2639 4573 2648 4607
rect 2596 4564 2648 4573
rect 2964 4428 3016 4480
rect 3884 4428 3936 4480
rect 2523 4326 2575 4378
rect 2587 4326 2639 4378
rect 2651 4326 2703 4378
rect 2715 4326 2767 4378
rect 4065 4326 4117 4378
rect 4129 4326 4181 4378
rect 4193 4326 4245 4378
rect 4257 4326 4309 4378
rect 2872 4224 2924 4276
rect 4620 4224 4672 4276
rect 2136 4131 2188 4140
rect 2136 4097 2145 4131
rect 2145 4097 2179 4131
rect 2179 4097 2188 4131
rect 2136 4088 2188 4097
rect 2872 4088 2924 4140
rect 2228 4020 2280 4072
rect 4436 4088 4488 4140
rect 4528 4020 4580 4072
rect 1768 3952 1820 4004
rect 2504 3952 2556 4004
rect 2044 3884 2096 3936
rect 2320 3927 2372 3936
rect 2320 3893 2329 3927
rect 2329 3893 2363 3927
rect 2363 3893 2372 3927
rect 2320 3884 2372 3893
rect 1753 3782 1805 3834
rect 1817 3782 1869 3834
rect 1881 3782 1933 3834
rect 1945 3782 1997 3834
rect 3294 3782 3346 3834
rect 3358 3782 3410 3834
rect 3422 3782 3474 3834
rect 3486 3782 3538 3834
rect 4836 3782 4888 3834
rect 4900 3782 4952 3834
rect 4964 3782 5016 3834
rect 5028 3782 5080 3834
rect 1584 3723 1636 3732
rect 1584 3689 1593 3723
rect 1593 3689 1627 3723
rect 1627 3689 1636 3723
rect 1584 3680 1636 3689
rect 2136 3723 2188 3732
rect 2136 3689 2145 3723
rect 2145 3689 2179 3723
rect 2179 3689 2188 3723
rect 2136 3680 2188 3689
rect 2228 3680 2280 3732
rect 2504 3680 2556 3732
rect 3884 3723 3936 3732
rect 3884 3689 3893 3723
rect 3893 3689 3927 3723
rect 3927 3689 3936 3723
rect 3884 3680 3936 3689
rect 2412 3587 2464 3596
rect 2412 3553 2421 3587
rect 2421 3553 2455 3587
rect 2455 3553 2464 3587
rect 2412 3544 2464 3553
rect 2872 3476 2924 3528
rect 2523 3238 2575 3290
rect 2587 3238 2639 3290
rect 2651 3238 2703 3290
rect 2715 3238 2767 3290
rect 4065 3238 4117 3290
rect 4129 3238 4181 3290
rect 4193 3238 4245 3290
rect 4257 3238 4309 3290
rect 2044 3136 2096 3188
rect 2320 3136 2372 3188
rect 3792 3136 3844 3188
rect 4712 3068 4764 3120
rect 1400 3043 1452 3052
rect 1400 3009 1409 3043
rect 1409 3009 1443 3043
rect 1443 3009 1452 3043
rect 1400 3000 1452 3009
rect 2044 3000 2096 3052
rect 2964 3000 3016 3052
rect 3148 3000 3200 3052
rect 3884 3000 3936 3052
rect 2872 2932 2924 2984
rect 4712 2796 4764 2848
rect 1753 2694 1805 2746
rect 1817 2694 1869 2746
rect 1881 2694 1933 2746
rect 1945 2694 1997 2746
rect 3294 2694 3346 2746
rect 3358 2694 3410 2746
rect 3422 2694 3474 2746
rect 3486 2694 3538 2746
rect 4836 2694 4888 2746
rect 4900 2694 4952 2746
rect 4964 2694 5016 2746
rect 5028 2694 5080 2746
rect 2872 2635 2924 2644
rect 2872 2601 2881 2635
rect 2881 2601 2915 2635
rect 2915 2601 2924 2635
rect 2872 2592 2924 2601
rect 3608 2592 3660 2644
rect 4436 2592 4488 2644
rect 2228 2456 2280 2508
rect 20 2388 72 2440
rect 2044 2388 2096 2440
rect 4068 2431 4120 2440
rect 4068 2397 4077 2431
rect 4077 2397 4111 2431
rect 4111 2397 4120 2431
rect 4068 2388 4120 2397
rect 4712 2388 4764 2440
rect 6092 2320 6144 2372
rect 2523 2150 2575 2202
rect 2587 2150 2639 2202
rect 2651 2150 2703 2202
rect 2715 2150 2767 2202
rect 4065 2150 4117 2202
rect 4129 2150 4181 2202
rect 4193 2150 4245 2202
rect 4257 2150 4309 2202
<< metal2 >>
rect 570 10177 626 10977
rect 2240 10254 2544 10282
rect 584 8566 612 10177
rect 1490 8800 1546 8809
rect 1490 8735 1546 8744
rect 1504 8634 1532 8735
rect 1492 8628 1544 8634
rect 1492 8570 1544 8576
rect 572 8560 624 8566
rect 572 8502 624 8508
rect 1584 8492 1636 8498
rect 1584 8434 1636 8440
rect 1596 8090 1624 8434
rect 1727 8188 2023 8208
rect 1783 8186 1807 8188
rect 1863 8186 1887 8188
rect 1943 8186 1967 8188
rect 1805 8134 1807 8186
rect 1869 8134 1881 8186
rect 1943 8134 1945 8186
rect 1783 8132 1807 8134
rect 1863 8132 1887 8134
rect 1943 8132 1967 8134
rect 1727 8112 2023 8132
rect 1584 8084 1636 8090
rect 1584 8026 1636 8032
rect 1492 7812 1544 7818
rect 1492 7754 1544 7760
rect 1504 7342 1532 7754
rect 2240 7426 2268 10254
rect 2516 10146 2544 10254
rect 2594 10177 2650 10977
rect 4618 10177 4674 10977
rect 6642 10177 6698 10977
rect 2608 10146 2636 10177
rect 2516 10118 2636 10146
rect 2497 8732 2793 8752
rect 2553 8730 2577 8732
rect 2633 8730 2657 8732
rect 2713 8730 2737 8732
rect 2575 8678 2577 8730
rect 2639 8678 2651 8730
rect 2713 8678 2715 8730
rect 2553 8676 2577 8678
rect 2633 8676 2657 8678
rect 2713 8676 2737 8678
rect 2497 8656 2793 8676
rect 4039 8732 4335 8752
rect 4095 8730 4119 8732
rect 4175 8730 4199 8732
rect 4255 8730 4279 8732
rect 4117 8678 4119 8730
rect 4181 8678 4193 8730
rect 4255 8678 4257 8730
rect 4095 8676 4119 8678
rect 4175 8676 4199 8678
rect 4255 8676 4279 8678
rect 4039 8656 4335 8676
rect 2320 8492 2372 8498
rect 2320 8434 2372 8440
rect 3884 8492 3936 8498
rect 3884 8434 3936 8440
rect 2332 7546 2360 8434
rect 3608 8288 3660 8294
rect 3608 8230 3660 8236
rect 3268 8188 3564 8208
rect 3324 8186 3348 8188
rect 3404 8186 3428 8188
rect 3484 8186 3508 8188
rect 3346 8134 3348 8186
rect 3410 8134 3422 8186
rect 3484 8134 3486 8186
rect 3324 8132 3348 8134
rect 3404 8132 3428 8134
rect 3484 8132 3508 8134
rect 3268 8112 3564 8132
rect 2412 7880 2464 7886
rect 2412 7822 2464 7828
rect 2320 7540 2372 7546
rect 2320 7482 2372 7488
rect 2136 7404 2188 7410
rect 2240 7398 2360 7426
rect 2136 7346 2188 7352
rect 1492 7336 1544 7342
rect 1492 7278 1544 7284
rect 1504 6914 1532 7278
rect 1727 7100 2023 7120
rect 1783 7098 1807 7100
rect 1863 7098 1887 7100
rect 1943 7098 1967 7100
rect 1805 7046 1807 7098
rect 1869 7046 1881 7098
rect 1943 7046 1945 7098
rect 1783 7044 1807 7046
rect 1863 7044 1887 7046
rect 1943 7044 1967 7046
rect 1727 7024 2023 7044
rect 1584 6928 1636 6934
rect 1504 6886 1584 6914
rect 1584 6870 1636 6876
rect 1400 6792 1452 6798
rect 1400 6734 1452 6740
rect 1412 5817 1440 6734
rect 1492 6656 1544 6662
rect 1492 6598 1544 6604
rect 1398 5808 1454 5817
rect 1398 5743 1454 5752
rect 1400 5704 1452 5710
rect 1400 5646 1452 5652
rect 1412 4826 1440 5646
rect 1504 5234 1532 6598
rect 1596 5778 1624 6870
rect 2044 6724 2096 6730
rect 2044 6666 2096 6672
rect 2056 6186 2084 6666
rect 2148 6390 2176 7346
rect 2228 6860 2280 6866
rect 2228 6802 2280 6808
rect 2136 6384 2188 6390
rect 2136 6326 2188 6332
rect 2044 6180 2096 6186
rect 2044 6122 2096 6128
rect 1727 6012 2023 6032
rect 1783 6010 1807 6012
rect 1863 6010 1887 6012
rect 1943 6010 1967 6012
rect 1805 5958 1807 6010
rect 1869 5958 1881 6010
rect 1943 5958 1945 6010
rect 1783 5956 1807 5958
rect 1863 5956 1887 5958
rect 1943 5956 1967 5958
rect 1727 5936 2023 5956
rect 1584 5772 1636 5778
rect 1584 5714 1636 5720
rect 2056 5710 2084 6122
rect 2044 5704 2096 5710
rect 2044 5646 2096 5652
rect 1492 5228 1544 5234
rect 1492 5170 1544 5176
rect 2136 5228 2188 5234
rect 2136 5170 2188 5176
rect 1727 4924 2023 4944
rect 1783 4922 1807 4924
rect 1863 4922 1887 4924
rect 1943 4922 1967 4924
rect 1805 4870 1807 4922
rect 1869 4870 1881 4922
rect 1943 4870 1945 4922
rect 1783 4868 1807 4870
rect 1863 4868 1887 4870
rect 1943 4868 1967 4870
rect 1727 4848 2023 4868
rect 1400 4820 1452 4826
rect 1400 4762 1452 4768
rect 2148 4622 2176 5170
rect 1584 4616 1636 4622
rect 1584 4558 1636 4564
rect 1768 4616 1820 4622
rect 1768 4558 1820 4564
rect 2136 4616 2188 4622
rect 2136 4558 2188 4564
rect 1596 3738 1624 4558
rect 1780 4010 1808 4558
rect 2148 4298 2176 4558
rect 2056 4270 2176 4298
rect 1768 4004 1820 4010
rect 1768 3946 1820 3952
rect 2056 3942 2084 4270
rect 2136 4140 2188 4146
rect 2136 4082 2188 4088
rect 2044 3936 2096 3942
rect 2044 3878 2096 3884
rect 1727 3836 2023 3856
rect 1783 3834 1807 3836
rect 1863 3834 1887 3836
rect 1943 3834 1967 3836
rect 1805 3782 1807 3834
rect 1869 3782 1881 3834
rect 1943 3782 1945 3834
rect 1783 3780 1807 3782
rect 1863 3780 1887 3782
rect 1943 3780 1967 3782
rect 1727 3760 2023 3780
rect 1584 3732 1636 3738
rect 1584 3674 1636 3680
rect 2056 3194 2084 3878
rect 2148 3738 2176 4082
rect 2240 4078 2268 6802
rect 2332 5642 2360 7398
rect 2424 7002 2452 7822
rect 3620 7818 3648 8230
rect 3896 7886 3924 8434
rect 4068 8356 4120 8362
rect 4068 8298 4120 8304
rect 4080 7886 4108 8298
rect 4436 8016 4488 8022
rect 4436 7958 4488 7964
rect 3884 7880 3936 7886
rect 3884 7822 3936 7828
rect 4068 7880 4120 7886
rect 4068 7822 4120 7828
rect 3608 7812 3660 7818
rect 3608 7754 3660 7760
rect 2497 7644 2793 7664
rect 2553 7642 2577 7644
rect 2633 7642 2657 7644
rect 2713 7642 2737 7644
rect 2575 7590 2577 7642
rect 2639 7590 2651 7642
rect 2713 7590 2715 7642
rect 2553 7588 2577 7590
rect 2633 7588 2657 7590
rect 2713 7588 2737 7590
rect 2497 7568 2793 7588
rect 3620 7410 3648 7754
rect 3792 7744 3844 7750
rect 3792 7686 3844 7692
rect 3608 7404 3660 7410
rect 3608 7346 3660 7352
rect 3608 7268 3660 7274
rect 3608 7210 3660 7216
rect 2780 7200 2832 7206
rect 2780 7142 2832 7148
rect 2412 6996 2464 7002
rect 2412 6938 2464 6944
rect 2792 6866 2820 7142
rect 3268 7100 3564 7120
rect 3324 7098 3348 7100
rect 3404 7098 3428 7100
rect 3484 7098 3508 7100
rect 3346 7046 3348 7098
rect 3410 7046 3422 7098
rect 3484 7046 3486 7098
rect 3324 7044 3348 7046
rect 3404 7044 3428 7046
rect 3484 7044 3508 7046
rect 3268 7024 3564 7044
rect 3620 7002 3648 7210
rect 3700 7200 3752 7206
rect 3700 7142 3752 7148
rect 3608 6996 3660 7002
rect 3608 6938 3660 6944
rect 2780 6860 2832 6866
rect 2780 6802 2832 6808
rect 3608 6860 3660 6866
rect 3608 6802 3660 6808
rect 2412 6792 2464 6798
rect 2412 6734 2464 6740
rect 3148 6792 3200 6798
rect 3148 6734 3200 6740
rect 2424 6322 2452 6734
rect 2872 6724 2924 6730
rect 2872 6666 2924 6672
rect 2497 6556 2793 6576
rect 2553 6554 2577 6556
rect 2633 6554 2657 6556
rect 2713 6554 2737 6556
rect 2575 6502 2577 6554
rect 2639 6502 2651 6554
rect 2713 6502 2715 6554
rect 2553 6500 2577 6502
rect 2633 6500 2657 6502
rect 2713 6500 2737 6502
rect 2497 6480 2793 6500
rect 2412 6316 2464 6322
rect 2412 6258 2464 6264
rect 2412 6180 2464 6186
rect 2412 6122 2464 6128
rect 2320 5636 2372 5642
rect 2320 5578 2372 5584
rect 2424 5574 2452 6122
rect 2884 5914 2912 6666
rect 2964 6656 3016 6662
rect 2964 6598 3016 6604
rect 2976 6390 3004 6598
rect 3160 6458 3188 6734
rect 3148 6452 3200 6458
rect 3148 6394 3200 6400
rect 2964 6384 3016 6390
rect 2964 6326 3016 6332
rect 3056 6316 3108 6322
rect 3056 6258 3108 6264
rect 2964 6248 3016 6254
rect 2964 6190 3016 6196
rect 2872 5908 2924 5914
rect 2872 5850 2924 5856
rect 2412 5568 2464 5574
rect 2412 5510 2464 5516
rect 2424 5370 2452 5510
rect 2497 5468 2793 5488
rect 2553 5466 2577 5468
rect 2633 5466 2657 5468
rect 2713 5466 2737 5468
rect 2575 5414 2577 5466
rect 2639 5414 2651 5466
rect 2713 5414 2715 5466
rect 2553 5412 2577 5414
rect 2633 5412 2657 5414
rect 2713 5412 2737 5414
rect 2497 5392 2793 5412
rect 2412 5364 2464 5370
rect 2412 5306 2464 5312
rect 2596 5296 2648 5302
rect 2596 5238 2648 5244
rect 2608 4622 2636 5238
rect 2780 5228 2832 5234
rect 2780 5170 2832 5176
rect 2792 4826 2820 5170
rect 2780 4820 2832 4826
rect 2780 4762 2832 4768
rect 2976 4758 3004 6190
rect 3068 5370 3096 6258
rect 3160 5710 3188 6394
rect 3268 6012 3564 6032
rect 3324 6010 3348 6012
rect 3404 6010 3428 6012
rect 3484 6010 3508 6012
rect 3346 5958 3348 6010
rect 3410 5958 3422 6010
rect 3484 5958 3486 6010
rect 3324 5956 3348 5958
rect 3404 5956 3428 5958
rect 3484 5956 3508 5958
rect 3268 5936 3564 5956
rect 3148 5704 3200 5710
rect 3148 5646 3200 5652
rect 3148 5568 3200 5574
rect 3148 5510 3200 5516
rect 3056 5364 3108 5370
rect 3056 5306 3108 5312
rect 3056 5160 3108 5166
rect 3056 5102 3108 5108
rect 2964 4752 3016 4758
rect 2964 4694 3016 4700
rect 2872 4684 2924 4690
rect 2872 4626 2924 4632
rect 2596 4616 2648 4622
rect 2424 4564 2596 4570
rect 2424 4558 2648 4564
rect 2424 4542 2636 4558
rect 2228 4072 2280 4078
rect 2228 4014 2280 4020
rect 2320 3936 2372 3942
rect 2320 3878 2372 3884
rect 2136 3732 2188 3738
rect 2136 3674 2188 3680
rect 2228 3732 2280 3738
rect 2228 3674 2280 3680
rect 2044 3188 2096 3194
rect 2044 3130 2096 3136
rect 2056 3058 2084 3130
rect 1400 3052 1452 3058
rect 1400 2994 1452 3000
rect 2044 3052 2096 3058
rect 2044 2994 2096 3000
rect 1412 2825 1440 2994
rect 1398 2816 1454 2825
rect 1398 2751 1454 2760
rect 1727 2748 2023 2768
rect 1783 2746 1807 2748
rect 1863 2746 1887 2748
rect 1943 2746 1967 2748
rect 1805 2694 1807 2746
rect 1869 2694 1881 2746
rect 1943 2694 1945 2746
rect 1783 2692 1807 2694
rect 1863 2692 1887 2694
rect 1943 2692 1967 2694
rect 1727 2672 2023 2692
rect 2240 2514 2268 3674
rect 2332 3194 2360 3878
rect 2424 3602 2452 4542
rect 2497 4380 2793 4400
rect 2553 4378 2577 4380
rect 2633 4378 2657 4380
rect 2713 4378 2737 4380
rect 2575 4326 2577 4378
rect 2639 4326 2651 4378
rect 2713 4326 2715 4378
rect 2553 4324 2577 4326
rect 2633 4324 2657 4326
rect 2713 4324 2737 4326
rect 2497 4304 2793 4324
rect 2884 4282 2912 4626
rect 3068 4570 3096 5102
rect 2976 4542 3096 4570
rect 2976 4486 3004 4542
rect 2964 4480 3016 4486
rect 2964 4422 3016 4428
rect 2872 4276 2924 4282
rect 2872 4218 2924 4224
rect 2884 4146 2912 4218
rect 2872 4140 2924 4146
rect 2872 4082 2924 4088
rect 2504 4004 2556 4010
rect 2504 3946 2556 3952
rect 2516 3738 2544 3946
rect 2504 3732 2556 3738
rect 2504 3674 2556 3680
rect 2412 3596 2464 3602
rect 2412 3538 2464 3544
rect 2884 3534 2912 4082
rect 2872 3528 2924 3534
rect 2872 3470 2924 3476
rect 2497 3292 2793 3312
rect 2553 3290 2577 3292
rect 2633 3290 2657 3292
rect 2713 3290 2737 3292
rect 2575 3238 2577 3290
rect 2639 3238 2651 3290
rect 2713 3238 2715 3290
rect 2553 3236 2577 3238
rect 2633 3236 2657 3238
rect 2713 3236 2737 3238
rect 2497 3216 2793 3236
rect 2320 3188 2372 3194
rect 2320 3130 2372 3136
rect 2976 3058 3004 4422
rect 3160 3058 3188 5510
rect 3268 4924 3564 4944
rect 3324 4922 3348 4924
rect 3404 4922 3428 4924
rect 3484 4922 3508 4924
rect 3346 4870 3348 4922
rect 3410 4870 3422 4922
rect 3484 4870 3486 4922
rect 3324 4868 3348 4870
rect 3404 4868 3428 4870
rect 3484 4868 3508 4870
rect 3268 4848 3564 4868
rect 3268 3836 3564 3856
rect 3324 3834 3348 3836
rect 3404 3834 3428 3836
rect 3484 3834 3508 3836
rect 3346 3782 3348 3834
rect 3410 3782 3422 3834
rect 3484 3782 3486 3834
rect 3324 3780 3348 3782
rect 3404 3780 3428 3782
rect 3484 3780 3508 3782
rect 3268 3760 3564 3780
rect 2964 3052 3016 3058
rect 2964 2994 3016 3000
rect 3148 3052 3200 3058
rect 3148 2994 3200 3000
rect 2872 2984 2924 2990
rect 2872 2926 2924 2932
rect 2884 2650 2912 2926
rect 3268 2748 3564 2768
rect 3324 2746 3348 2748
rect 3404 2746 3428 2748
rect 3484 2746 3508 2748
rect 3346 2694 3348 2746
rect 3410 2694 3422 2746
rect 3484 2694 3486 2746
rect 3324 2692 3348 2694
rect 3404 2692 3428 2694
rect 3484 2692 3508 2694
rect 3268 2672 3564 2692
rect 3620 2650 3648 6802
rect 3712 6390 3740 7142
rect 3804 6934 3832 7686
rect 3896 7410 3924 7822
rect 4039 7644 4335 7664
rect 4095 7642 4119 7644
rect 4175 7642 4199 7644
rect 4255 7642 4279 7644
rect 4117 7590 4119 7642
rect 4181 7590 4193 7642
rect 4255 7590 4257 7642
rect 4095 7588 4119 7590
rect 4175 7588 4199 7590
rect 4255 7588 4279 7590
rect 4039 7568 4335 7588
rect 3884 7404 3936 7410
rect 3884 7346 3936 7352
rect 3792 6928 3844 6934
rect 3792 6870 3844 6876
rect 3700 6384 3752 6390
rect 3700 6326 3752 6332
rect 3712 5030 3740 6326
rect 3896 6254 3924 7346
rect 4448 7206 4476 7958
rect 4528 7336 4580 7342
rect 4528 7278 4580 7284
rect 4436 7200 4488 7206
rect 4436 7142 4488 7148
rect 4540 7018 4568 7278
rect 4448 7002 4568 7018
rect 4436 6996 4568 7002
rect 4488 6990 4568 6996
rect 4436 6938 4488 6944
rect 4039 6556 4335 6576
rect 4095 6554 4119 6556
rect 4175 6554 4199 6556
rect 4255 6554 4279 6556
rect 4117 6502 4119 6554
rect 4181 6502 4193 6554
rect 4255 6502 4257 6554
rect 4095 6500 4119 6502
rect 4175 6500 4199 6502
rect 4255 6500 4279 6502
rect 4039 6480 4335 6500
rect 3976 6316 4028 6322
rect 3976 6258 4028 6264
rect 3884 6248 3936 6254
rect 3884 6190 3936 6196
rect 3792 5568 3844 5574
rect 3792 5510 3844 5516
rect 3804 5234 3832 5510
rect 3792 5228 3844 5234
rect 3792 5170 3844 5176
rect 3896 5166 3924 6190
rect 3988 5778 4016 6258
rect 4448 6118 4476 6938
rect 4632 6798 4660 10177
rect 4712 8424 4764 8430
rect 4712 8366 4764 8372
rect 4724 7886 4752 8366
rect 5540 8288 5592 8294
rect 5540 8230 5592 8236
rect 4810 8188 5106 8208
rect 4866 8186 4890 8188
rect 4946 8186 4970 8188
rect 5026 8186 5050 8188
rect 4888 8134 4890 8186
rect 4952 8134 4964 8186
rect 5026 8134 5028 8186
rect 4866 8132 4890 8134
rect 4946 8132 4970 8134
rect 5026 8132 5050 8134
rect 4810 8112 5106 8132
rect 5552 7993 5580 8230
rect 5538 7984 5594 7993
rect 5538 7919 5594 7928
rect 4712 7880 4764 7886
rect 4712 7822 4764 7828
rect 4712 7268 4764 7274
rect 4712 7210 4764 7216
rect 4724 6866 4752 7210
rect 4810 7100 5106 7120
rect 4866 7098 4890 7100
rect 4946 7098 4970 7100
rect 5026 7098 5050 7100
rect 4888 7046 4890 7098
rect 4952 7046 4964 7098
rect 5026 7046 5028 7098
rect 4866 7044 4890 7046
rect 4946 7044 4970 7046
rect 5026 7044 5050 7046
rect 4810 7024 5106 7044
rect 4712 6860 4764 6866
rect 4712 6802 4764 6808
rect 4620 6792 4672 6798
rect 4620 6734 4672 6740
rect 4528 6656 4580 6662
rect 4528 6598 4580 6604
rect 4436 6112 4488 6118
rect 4436 6054 4488 6060
rect 3976 5772 4028 5778
rect 3976 5714 4028 5720
rect 4436 5772 4488 5778
rect 4436 5714 4488 5720
rect 4039 5468 4335 5488
rect 4095 5466 4119 5468
rect 4175 5466 4199 5468
rect 4255 5466 4279 5468
rect 4117 5414 4119 5466
rect 4181 5414 4193 5466
rect 4255 5414 4257 5466
rect 4095 5412 4119 5414
rect 4175 5412 4199 5414
rect 4255 5412 4279 5414
rect 4039 5392 4335 5412
rect 3884 5160 3936 5166
rect 3804 5108 3884 5114
rect 3804 5102 3936 5108
rect 3804 5086 3924 5102
rect 3700 5024 3752 5030
rect 3700 4966 3752 4972
rect 3804 3194 3832 5086
rect 3884 4480 3936 4486
rect 3884 4422 3936 4428
rect 3896 3738 3924 4422
rect 4039 4380 4335 4400
rect 4095 4378 4119 4380
rect 4175 4378 4199 4380
rect 4255 4378 4279 4380
rect 4117 4326 4119 4378
rect 4181 4326 4193 4378
rect 4255 4326 4257 4378
rect 4095 4324 4119 4326
rect 4175 4324 4199 4326
rect 4255 4324 4279 4326
rect 4039 4304 4335 4324
rect 4448 4146 4476 5714
rect 4540 4690 4568 6598
rect 4724 6458 4752 6802
rect 4712 6452 4764 6458
rect 4712 6394 4764 6400
rect 4712 6316 4764 6322
rect 4712 6258 4764 6264
rect 4620 6112 4672 6118
rect 4620 6054 4672 6060
rect 4632 5710 4660 6054
rect 4620 5704 4672 5710
rect 4620 5646 4672 5652
rect 4528 4684 4580 4690
rect 4528 4626 4580 4632
rect 4436 4140 4488 4146
rect 4436 4082 4488 4088
rect 3884 3732 3936 3738
rect 3884 3674 3936 3680
rect 4039 3292 4335 3312
rect 4095 3290 4119 3292
rect 4175 3290 4199 3292
rect 4255 3290 4279 3292
rect 4117 3238 4119 3290
rect 4181 3238 4193 3290
rect 4255 3238 4257 3290
rect 4095 3236 4119 3238
rect 4175 3236 4199 3238
rect 4255 3236 4279 3238
rect 4039 3216 4335 3236
rect 3792 3188 3844 3194
rect 3792 3130 3844 3136
rect 3884 3052 3936 3058
rect 3884 2994 3936 3000
rect 2872 2644 2924 2650
rect 2872 2586 2924 2592
rect 3608 2644 3660 2650
rect 3608 2586 3660 2592
rect 2228 2508 2280 2514
rect 2228 2450 2280 2456
rect 20 2440 72 2446
rect 20 2382 72 2388
rect 2044 2440 2096 2446
rect 2044 2382 2096 2388
rect 32 800 60 2382
rect 2056 800 2084 2382
rect 2497 2204 2793 2224
rect 2553 2202 2577 2204
rect 2633 2202 2657 2204
rect 2713 2202 2737 2204
rect 2575 2150 2577 2202
rect 2639 2150 2651 2202
rect 2713 2150 2715 2202
rect 2553 2148 2577 2150
rect 2633 2148 2657 2150
rect 2713 2148 2737 2150
rect 2497 2128 2793 2148
rect 3896 1578 3924 2994
rect 4448 2650 4476 4082
rect 4540 4078 4568 4626
rect 4632 4282 4660 5646
rect 4724 5642 4752 6258
rect 4810 6012 5106 6032
rect 4866 6010 4890 6012
rect 4946 6010 4970 6012
rect 5026 6010 5050 6012
rect 4888 5958 4890 6010
rect 4952 5958 4964 6010
rect 5026 5958 5028 6010
rect 4866 5956 4890 5958
rect 4946 5956 4970 5958
rect 5026 5956 5050 5958
rect 4810 5936 5106 5956
rect 6656 5846 6684 10177
rect 6644 5840 6696 5846
rect 6644 5782 6696 5788
rect 4712 5636 4764 5642
rect 4712 5578 4764 5584
rect 4620 4276 4672 4282
rect 4620 4218 4672 4224
rect 4528 4072 4580 4078
rect 4528 4014 4580 4020
rect 4724 3126 4752 5578
rect 4804 5568 4856 5574
rect 4804 5510 4856 5516
rect 4816 5302 4844 5510
rect 4804 5296 4856 5302
rect 4804 5238 4856 5244
rect 5356 5092 5408 5098
rect 5356 5034 5408 5040
rect 5368 5001 5396 5034
rect 5354 4992 5410 5001
rect 4810 4924 5106 4944
rect 5354 4927 5410 4936
rect 4866 4922 4890 4924
rect 4946 4922 4970 4924
rect 5026 4922 5050 4924
rect 4888 4870 4890 4922
rect 4952 4870 4964 4922
rect 5026 4870 5028 4922
rect 4866 4868 4890 4870
rect 4946 4868 4970 4870
rect 5026 4868 5050 4870
rect 4810 4848 5106 4868
rect 4810 3836 5106 3856
rect 4866 3834 4890 3836
rect 4946 3834 4970 3836
rect 5026 3834 5050 3836
rect 4888 3782 4890 3834
rect 4952 3782 4964 3834
rect 5026 3782 5028 3834
rect 4866 3780 4890 3782
rect 4946 3780 4970 3782
rect 5026 3780 5050 3782
rect 4810 3760 5106 3780
rect 4712 3120 4764 3126
rect 4712 3062 4764 3068
rect 4712 2848 4764 2854
rect 4712 2790 4764 2796
rect 4436 2644 4488 2650
rect 4436 2586 4488 2592
rect 4724 2446 4752 2790
rect 4810 2748 5106 2768
rect 4866 2746 4890 2748
rect 4946 2746 4970 2748
rect 5026 2746 5050 2748
rect 4888 2694 4890 2746
rect 4952 2694 4964 2746
rect 5026 2694 5028 2746
rect 4866 2692 4890 2694
rect 4946 2692 4970 2694
rect 5026 2692 5050 2694
rect 4810 2672 5106 2692
rect 4068 2440 4120 2446
rect 4066 2408 4068 2417
rect 4712 2440 4764 2446
rect 4120 2408 4122 2417
rect 4712 2382 4764 2388
rect 4066 2343 4122 2352
rect 6092 2372 6144 2378
rect 6092 2314 6144 2320
rect 4039 2204 4335 2224
rect 4095 2202 4119 2204
rect 4175 2202 4199 2204
rect 4255 2202 4279 2204
rect 4117 2150 4119 2202
rect 4181 2150 4193 2202
rect 4255 2150 4257 2202
rect 4095 2148 4119 2150
rect 4175 2148 4199 2150
rect 4255 2148 4279 2150
rect 4039 2128 4335 2148
rect 3896 1550 4108 1578
rect 4080 800 4108 1550
rect 6104 800 6132 2314
rect 18 0 74 800
rect 2042 0 2098 800
rect 4066 0 4122 800
rect 6090 0 6146 800
<< via2 >>
rect 1490 8744 1546 8800
rect 1727 8186 1783 8188
rect 1807 8186 1863 8188
rect 1887 8186 1943 8188
rect 1967 8186 2023 8188
rect 1727 8134 1753 8186
rect 1753 8134 1783 8186
rect 1807 8134 1817 8186
rect 1817 8134 1863 8186
rect 1887 8134 1933 8186
rect 1933 8134 1943 8186
rect 1967 8134 1997 8186
rect 1997 8134 2023 8186
rect 1727 8132 1783 8134
rect 1807 8132 1863 8134
rect 1887 8132 1943 8134
rect 1967 8132 2023 8134
rect 2497 8730 2553 8732
rect 2577 8730 2633 8732
rect 2657 8730 2713 8732
rect 2737 8730 2793 8732
rect 2497 8678 2523 8730
rect 2523 8678 2553 8730
rect 2577 8678 2587 8730
rect 2587 8678 2633 8730
rect 2657 8678 2703 8730
rect 2703 8678 2713 8730
rect 2737 8678 2767 8730
rect 2767 8678 2793 8730
rect 2497 8676 2553 8678
rect 2577 8676 2633 8678
rect 2657 8676 2713 8678
rect 2737 8676 2793 8678
rect 4039 8730 4095 8732
rect 4119 8730 4175 8732
rect 4199 8730 4255 8732
rect 4279 8730 4335 8732
rect 4039 8678 4065 8730
rect 4065 8678 4095 8730
rect 4119 8678 4129 8730
rect 4129 8678 4175 8730
rect 4199 8678 4245 8730
rect 4245 8678 4255 8730
rect 4279 8678 4309 8730
rect 4309 8678 4335 8730
rect 4039 8676 4095 8678
rect 4119 8676 4175 8678
rect 4199 8676 4255 8678
rect 4279 8676 4335 8678
rect 3268 8186 3324 8188
rect 3348 8186 3404 8188
rect 3428 8186 3484 8188
rect 3508 8186 3564 8188
rect 3268 8134 3294 8186
rect 3294 8134 3324 8186
rect 3348 8134 3358 8186
rect 3358 8134 3404 8186
rect 3428 8134 3474 8186
rect 3474 8134 3484 8186
rect 3508 8134 3538 8186
rect 3538 8134 3564 8186
rect 3268 8132 3324 8134
rect 3348 8132 3404 8134
rect 3428 8132 3484 8134
rect 3508 8132 3564 8134
rect 1727 7098 1783 7100
rect 1807 7098 1863 7100
rect 1887 7098 1943 7100
rect 1967 7098 2023 7100
rect 1727 7046 1753 7098
rect 1753 7046 1783 7098
rect 1807 7046 1817 7098
rect 1817 7046 1863 7098
rect 1887 7046 1933 7098
rect 1933 7046 1943 7098
rect 1967 7046 1997 7098
rect 1997 7046 2023 7098
rect 1727 7044 1783 7046
rect 1807 7044 1863 7046
rect 1887 7044 1943 7046
rect 1967 7044 2023 7046
rect 1398 5752 1454 5808
rect 1727 6010 1783 6012
rect 1807 6010 1863 6012
rect 1887 6010 1943 6012
rect 1967 6010 2023 6012
rect 1727 5958 1753 6010
rect 1753 5958 1783 6010
rect 1807 5958 1817 6010
rect 1817 5958 1863 6010
rect 1887 5958 1933 6010
rect 1933 5958 1943 6010
rect 1967 5958 1997 6010
rect 1997 5958 2023 6010
rect 1727 5956 1783 5958
rect 1807 5956 1863 5958
rect 1887 5956 1943 5958
rect 1967 5956 2023 5958
rect 1727 4922 1783 4924
rect 1807 4922 1863 4924
rect 1887 4922 1943 4924
rect 1967 4922 2023 4924
rect 1727 4870 1753 4922
rect 1753 4870 1783 4922
rect 1807 4870 1817 4922
rect 1817 4870 1863 4922
rect 1887 4870 1933 4922
rect 1933 4870 1943 4922
rect 1967 4870 1997 4922
rect 1997 4870 2023 4922
rect 1727 4868 1783 4870
rect 1807 4868 1863 4870
rect 1887 4868 1943 4870
rect 1967 4868 2023 4870
rect 1727 3834 1783 3836
rect 1807 3834 1863 3836
rect 1887 3834 1943 3836
rect 1967 3834 2023 3836
rect 1727 3782 1753 3834
rect 1753 3782 1783 3834
rect 1807 3782 1817 3834
rect 1817 3782 1863 3834
rect 1887 3782 1933 3834
rect 1933 3782 1943 3834
rect 1967 3782 1997 3834
rect 1997 3782 2023 3834
rect 1727 3780 1783 3782
rect 1807 3780 1863 3782
rect 1887 3780 1943 3782
rect 1967 3780 2023 3782
rect 2497 7642 2553 7644
rect 2577 7642 2633 7644
rect 2657 7642 2713 7644
rect 2737 7642 2793 7644
rect 2497 7590 2523 7642
rect 2523 7590 2553 7642
rect 2577 7590 2587 7642
rect 2587 7590 2633 7642
rect 2657 7590 2703 7642
rect 2703 7590 2713 7642
rect 2737 7590 2767 7642
rect 2767 7590 2793 7642
rect 2497 7588 2553 7590
rect 2577 7588 2633 7590
rect 2657 7588 2713 7590
rect 2737 7588 2793 7590
rect 3268 7098 3324 7100
rect 3348 7098 3404 7100
rect 3428 7098 3484 7100
rect 3508 7098 3564 7100
rect 3268 7046 3294 7098
rect 3294 7046 3324 7098
rect 3348 7046 3358 7098
rect 3358 7046 3404 7098
rect 3428 7046 3474 7098
rect 3474 7046 3484 7098
rect 3508 7046 3538 7098
rect 3538 7046 3564 7098
rect 3268 7044 3324 7046
rect 3348 7044 3404 7046
rect 3428 7044 3484 7046
rect 3508 7044 3564 7046
rect 2497 6554 2553 6556
rect 2577 6554 2633 6556
rect 2657 6554 2713 6556
rect 2737 6554 2793 6556
rect 2497 6502 2523 6554
rect 2523 6502 2553 6554
rect 2577 6502 2587 6554
rect 2587 6502 2633 6554
rect 2657 6502 2703 6554
rect 2703 6502 2713 6554
rect 2737 6502 2767 6554
rect 2767 6502 2793 6554
rect 2497 6500 2553 6502
rect 2577 6500 2633 6502
rect 2657 6500 2713 6502
rect 2737 6500 2793 6502
rect 2497 5466 2553 5468
rect 2577 5466 2633 5468
rect 2657 5466 2713 5468
rect 2737 5466 2793 5468
rect 2497 5414 2523 5466
rect 2523 5414 2553 5466
rect 2577 5414 2587 5466
rect 2587 5414 2633 5466
rect 2657 5414 2703 5466
rect 2703 5414 2713 5466
rect 2737 5414 2767 5466
rect 2767 5414 2793 5466
rect 2497 5412 2553 5414
rect 2577 5412 2633 5414
rect 2657 5412 2713 5414
rect 2737 5412 2793 5414
rect 3268 6010 3324 6012
rect 3348 6010 3404 6012
rect 3428 6010 3484 6012
rect 3508 6010 3564 6012
rect 3268 5958 3294 6010
rect 3294 5958 3324 6010
rect 3348 5958 3358 6010
rect 3358 5958 3404 6010
rect 3428 5958 3474 6010
rect 3474 5958 3484 6010
rect 3508 5958 3538 6010
rect 3538 5958 3564 6010
rect 3268 5956 3324 5958
rect 3348 5956 3404 5958
rect 3428 5956 3484 5958
rect 3508 5956 3564 5958
rect 1398 2760 1454 2816
rect 1727 2746 1783 2748
rect 1807 2746 1863 2748
rect 1887 2746 1943 2748
rect 1967 2746 2023 2748
rect 1727 2694 1753 2746
rect 1753 2694 1783 2746
rect 1807 2694 1817 2746
rect 1817 2694 1863 2746
rect 1887 2694 1933 2746
rect 1933 2694 1943 2746
rect 1967 2694 1997 2746
rect 1997 2694 2023 2746
rect 1727 2692 1783 2694
rect 1807 2692 1863 2694
rect 1887 2692 1943 2694
rect 1967 2692 2023 2694
rect 2497 4378 2553 4380
rect 2577 4378 2633 4380
rect 2657 4378 2713 4380
rect 2737 4378 2793 4380
rect 2497 4326 2523 4378
rect 2523 4326 2553 4378
rect 2577 4326 2587 4378
rect 2587 4326 2633 4378
rect 2657 4326 2703 4378
rect 2703 4326 2713 4378
rect 2737 4326 2767 4378
rect 2767 4326 2793 4378
rect 2497 4324 2553 4326
rect 2577 4324 2633 4326
rect 2657 4324 2713 4326
rect 2737 4324 2793 4326
rect 2497 3290 2553 3292
rect 2577 3290 2633 3292
rect 2657 3290 2713 3292
rect 2737 3290 2793 3292
rect 2497 3238 2523 3290
rect 2523 3238 2553 3290
rect 2577 3238 2587 3290
rect 2587 3238 2633 3290
rect 2657 3238 2703 3290
rect 2703 3238 2713 3290
rect 2737 3238 2767 3290
rect 2767 3238 2793 3290
rect 2497 3236 2553 3238
rect 2577 3236 2633 3238
rect 2657 3236 2713 3238
rect 2737 3236 2793 3238
rect 3268 4922 3324 4924
rect 3348 4922 3404 4924
rect 3428 4922 3484 4924
rect 3508 4922 3564 4924
rect 3268 4870 3294 4922
rect 3294 4870 3324 4922
rect 3348 4870 3358 4922
rect 3358 4870 3404 4922
rect 3428 4870 3474 4922
rect 3474 4870 3484 4922
rect 3508 4870 3538 4922
rect 3538 4870 3564 4922
rect 3268 4868 3324 4870
rect 3348 4868 3404 4870
rect 3428 4868 3484 4870
rect 3508 4868 3564 4870
rect 3268 3834 3324 3836
rect 3348 3834 3404 3836
rect 3428 3834 3484 3836
rect 3508 3834 3564 3836
rect 3268 3782 3294 3834
rect 3294 3782 3324 3834
rect 3348 3782 3358 3834
rect 3358 3782 3404 3834
rect 3428 3782 3474 3834
rect 3474 3782 3484 3834
rect 3508 3782 3538 3834
rect 3538 3782 3564 3834
rect 3268 3780 3324 3782
rect 3348 3780 3404 3782
rect 3428 3780 3484 3782
rect 3508 3780 3564 3782
rect 3268 2746 3324 2748
rect 3348 2746 3404 2748
rect 3428 2746 3484 2748
rect 3508 2746 3564 2748
rect 3268 2694 3294 2746
rect 3294 2694 3324 2746
rect 3348 2694 3358 2746
rect 3358 2694 3404 2746
rect 3428 2694 3474 2746
rect 3474 2694 3484 2746
rect 3508 2694 3538 2746
rect 3538 2694 3564 2746
rect 3268 2692 3324 2694
rect 3348 2692 3404 2694
rect 3428 2692 3484 2694
rect 3508 2692 3564 2694
rect 4039 7642 4095 7644
rect 4119 7642 4175 7644
rect 4199 7642 4255 7644
rect 4279 7642 4335 7644
rect 4039 7590 4065 7642
rect 4065 7590 4095 7642
rect 4119 7590 4129 7642
rect 4129 7590 4175 7642
rect 4199 7590 4245 7642
rect 4245 7590 4255 7642
rect 4279 7590 4309 7642
rect 4309 7590 4335 7642
rect 4039 7588 4095 7590
rect 4119 7588 4175 7590
rect 4199 7588 4255 7590
rect 4279 7588 4335 7590
rect 4039 6554 4095 6556
rect 4119 6554 4175 6556
rect 4199 6554 4255 6556
rect 4279 6554 4335 6556
rect 4039 6502 4065 6554
rect 4065 6502 4095 6554
rect 4119 6502 4129 6554
rect 4129 6502 4175 6554
rect 4199 6502 4245 6554
rect 4245 6502 4255 6554
rect 4279 6502 4309 6554
rect 4309 6502 4335 6554
rect 4039 6500 4095 6502
rect 4119 6500 4175 6502
rect 4199 6500 4255 6502
rect 4279 6500 4335 6502
rect 4810 8186 4866 8188
rect 4890 8186 4946 8188
rect 4970 8186 5026 8188
rect 5050 8186 5106 8188
rect 4810 8134 4836 8186
rect 4836 8134 4866 8186
rect 4890 8134 4900 8186
rect 4900 8134 4946 8186
rect 4970 8134 5016 8186
rect 5016 8134 5026 8186
rect 5050 8134 5080 8186
rect 5080 8134 5106 8186
rect 4810 8132 4866 8134
rect 4890 8132 4946 8134
rect 4970 8132 5026 8134
rect 5050 8132 5106 8134
rect 5538 7928 5594 7984
rect 4810 7098 4866 7100
rect 4890 7098 4946 7100
rect 4970 7098 5026 7100
rect 5050 7098 5106 7100
rect 4810 7046 4836 7098
rect 4836 7046 4866 7098
rect 4890 7046 4900 7098
rect 4900 7046 4946 7098
rect 4970 7046 5016 7098
rect 5016 7046 5026 7098
rect 5050 7046 5080 7098
rect 5080 7046 5106 7098
rect 4810 7044 4866 7046
rect 4890 7044 4946 7046
rect 4970 7044 5026 7046
rect 5050 7044 5106 7046
rect 4039 5466 4095 5468
rect 4119 5466 4175 5468
rect 4199 5466 4255 5468
rect 4279 5466 4335 5468
rect 4039 5414 4065 5466
rect 4065 5414 4095 5466
rect 4119 5414 4129 5466
rect 4129 5414 4175 5466
rect 4199 5414 4245 5466
rect 4245 5414 4255 5466
rect 4279 5414 4309 5466
rect 4309 5414 4335 5466
rect 4039 5412 4095 5414
rect 4119 5412 4175 5414
rect 4199 5412 4255 5414
rect 4279 5412 4335 5414
rect 4039 4378 4095 4380
rect 4119 4378 4175 4380
rect 4199 4378 4255 4380
rect 4279 4378 4335 4380
rect 4039 4326 4065 4378
rect 4065 4326 4095 4378
rect 4119 4326 4129 4378
rect 4129 4326 4175 4378
rect 4199 4326 4245 4378
rect 4245 4326 4255 4378
rect 4279 4326 4309 4378
rect 4309 4326 4335 4378
rect 4039 4324 4095 4326
rect 4119 4324 4175 4326
rect 4199 4324 4255 4326
rect 4279 4324 4335 4326
rect 4039 3290 4095 3292
rect 4119 3290 4175 3292
rect 4199 3290 4255 3292
rect 4279 3290 4335 3292
rect 4039 3238 4065 3290
rect 4065 3238 4095 3290
rect 4119 3238 4129 3290
rect 4129 3238 4175 3290
rect 4199 3238 4245 3290
rect 4245 3238 4255 3290
rect 4279 3238 4309 3290
rect 4309 3238 4335 3290
rect 4039 3236 4095 3238
rect 4119 3236 4175 3238
rect 4199 3236 4255 3238
rect 4279 3236 4335 3238
rect 2497 2202 2553 2204
rect 2577 2202 2633 2204
rect 2657 2202 2713 2204
rect 2737 2202 2793 2204
rect 2497 2150 2523 2202
rect 2523 2150 2553 2202
rect 2577 2150 2587 2202
rect 2587 2150 2633 2202
rect 2657 2150 2703 2202
rect 2703 2150 2713 2202
rect 2737 2150 2767 2202
rect 2767 2150 2793 2202
rect 2497 2148 2553 2150
rect 2577 2148 2633 2150
rect 2657 2148 2713 2150
rect 2737 2148 2793 2150
rect 4810 6010 4866 6012
rect 4890 6010 4946 6012
rect 4970 6010 5026 6012
rect 5050 6010 5106 6012
rect 4810 5958 4836 6010
rect 4836 5958 4866 6010
rect 4890 5958 4900 6010
rect 4900 5958 4946 6010
rect 4970 5958 5016 6010
rect 5016 5958 5026 6010
rect 5050 5958 5080 6010
rect 5080 5958 5106 6010
rect 4810 5956 4866 5958
rect 4890 5956 4946 5958
rect 4970 5956 5026 5958
rect 5050 5956 5106 5958
rect 5354 4936 5410 4992
rect 4810 4922 4866 4924
rect 4890 4922 4946 4924
rect 4970 4922 5026 4924
rect 5050 4922 5106 4924
rect 4810 4870 4836 4922
rect 4836 4870 4866 4922
rect 4890 4870 4900 4922
rect 4900 4870 4946 4922
rect 4970 4870 5016 4922
rect 5016 4870 5026 4922
rect 5050 4870 5080 4922
rect 5080 4870 5106 4922
rect 4810 4868 4866 4870
rect 4890 4868 4946 4870
rect 4970 4868 5026 4870
rect 5050 4868 5106 4870
rect 4810 3834 4866 3836
rect 4890 3834 4946 3836
rect 4970 3834 5026 3836
rect 5050 3834 5106 3836
rect 4810 3782 4836 3834
rect 4836 3782 4866 3834
rect 4890 3782 4900 3834
rect 4900 3782 4946 3834
rect 4970 3782 5016 3834
rect 5016 3782 5026 3834
rect 5050 3782 5080 3834
rect 5080 3782 5106 3834
rect 4810 3780 4866 3782
rect 4890 3780 4946 3782
rect 4970 3780 5026 3782
rect 5050 3780 5106 3782
rect 4810 2746 4866 2748
rect 4890 2746 4946 2748
rect 4970 2746 5026 2748
rect 5050 2746 5106 2748
rect 4810 2694 4836 2746
rect 4836 2694 4866 2746
rect 4890 2694 4900 2746
rect 4900 2694 4946 2746
rect 4970 2694 5016 2746
rect 5016 2694 5026 2746
rect 5050 2694 5080 2746
rect 5080 2694 5106 2746
rect 4810 2692 4866 2694
rect 4890 2692 4946 2694
rect 4970 2692 5026 2694
rect 5050 2692 5106 2694
rect 4066 2388 4068 2408
rect 4068 2388 4120 2408
rect 4120 2388 4122 2408
rect 4066 2352 4122 2388
rect 4039 2202 4095 2204
rect 4119 2202 4175 2204
rect 4199 2202 4255 2204
rect 4279 2202 4335 2204
rect 4039 2150 4065 2202
rect 4065 2150 4095 2202
rect 4119 2150 4129 2202
rect 4129 2150 4175 2202
rect 4199 2150 4245 2202
rect 4245 2150 4255 2202
rect 4279 2150 4309 2202
rect 4309 2150 4335 2202
rect 4039 2148 4095 2150
rect 4119 2148 4175 2150
rect 4199 2148 4255 2150
rect 4279 2148 4335 2150
<< metal3 >>
rect 0 8802 800 8832
rect 1485 8802 1551 8805
rect 0 8800 1551 8802
rect 0 8744 1490 8800
rect 1546 8744 1551 8800
rect 0 8742 1551 8744
rect 0 8712 800 8742
rect 1485 8739 1551 8742
rect 2485 8736 2805 8737
rect 2485 8672 2493 8736
rect 2557 8672 2573 8736
rect 2637 8672 2653 8736
rect 2717 8672 2733 8736
rect 2797 8672 2805 8736
rect 2485 8671 2805 8672
rect 4027 8736 4347 8737
rect 4027 8672 4035 8736
rect 4099 8672 4115 8736
rect 4179 8672 4195 8736
rect 4259 8672 4275 8736
rect 4339 8672 4347 8736
rect 4027 8671 4347 8672
rect 1715 8192 2035 8193
rect 1715 8128 1723 8192
rect 1787 8128 1803 8192
rect 1867 8128 1883 8192
rect 1947 8128 1963 8192
rect 2027 8128 2035 8192
rect 1715 8127 2035 8128
rect 3256 8192 3576 8193
rect 3256 8128 3264 8192
rect 3328 8128 3344 8192
rect 3408 8128 3424 8192
rect 3488 8128 3504 8192
rect 3568 8128 3576 8192
rect 3256 8127 3576 8128
rect 4798 8192 5118 8193
rect 4798 8128 4806 8192
rect 4870 8128 4886 8192
rect 4950 8128 4966 8192
rect 5030 8128 5046 8192
rect 5110 8128 5118 8192
rect 4798 8127 5118 8128
rect 5533 7986 5599 7989
rect 6033 7986 6833 8016
rect 5533 7984 6833 7986
rect 5533 7928 5538 7984
rect 5594 7928 6833 7984
rect 5533 7926 6833 7928
rect 5533 7923 5599 7926
rect 6033 7896 6833 7926
rect 2485 7648 2805 7649
rect 2485 7584 2493 7648
rect 2557 7584 2573 7648
rect 2637 7584 2653 7648
rect 2717 7584 2733 7648
rect 2797 7584 2805 7648
rect 2485 7583 2805 7584
rect 4027 7648 4347 7649
rect 4027 7584 4035 7648
rect 4099 7584 4115 7648
rect 4179 7584 4195 7648
rect 4259 7584 4275 7648
rect 4339 7584 4347 7648
rect 4027 7583 4347 7584
rect 1715 7104 2035 7105
rect 1715 7040 1723 7104
rect 1787 7040 1803 7104
rect 1867 7040 1883 7104
rect 1947 7040 1963 7104
rect 2027 7040 2035 7104
rect 1715 7039 2035 7040
rect 3256 7104 3576 7105
rect 3256 7040 3264 7104
rect 3328 7040 3344 7104
rect 3408 7040 3424 7104
rect 3488 7040 3504 7104
rect 3568 7040 3576 7104
rect 3256 7039 3576 7040
rect 4798 7104 5118 7105
rect 4798 7040 4806 7104
rect 4870 7040 4886 7104
rect 4950 7040 4966 7104
rect 5030 7040 5046 7104
rect 5110 7040 5118 7104
rect 4798 7039 5118 7040
rect 2485 6560 2805 6561
rect 2485 6496 2493 6560
rect 2557 6496 2573 6560
rect 2637 6496 2653 6560
rect 2717 6496 2733 6560
rect 2797 6496 2805 6560
rect 2485 6495 2805 6496
rect 4027 6560 4347 6561
rect 4027 6496 4035 6560
rect 4099 6496 4115 6560
rect 4179 6496 4195 6560
rect 4259 6496 4275 6560
rect 4339 6496 4347 6560
rect 4027 6495 4347 6496
rect 1715 6016 2035 6017
rect 1715 5952 1723 6016
rect 1787 5952 1803 6016
rect 1867 5952 1883 6016
rect 1947 5952 1963 6016
rect 2027 5952 2035 6016
rect 1715 5951 2035 5952
rect 3256 6016 3576 6017
rect 3256 5952 3264 6016
rect 3328 5952 3344 6016
rect 3408 5952 3424 6016
rect 3488 5952 3504 6016
rect 3568 5952 3576 6016
rect 3256 5951 3576 5952
rect 4798 6016 5118 6017
rect 4798 5952 4806 6016
rect 4870 5952 4886 6016
rect 4950 5952 4966 6016
rect 5030 5952 5046 6016
rect 5110 5952 5118 6016
rect 4798 5951 5118 5952
rect 0 5810 800 5840
rect 1393 5810 1459 5813
rect 0 5808 1459 5810
rect 0 5752 1398 5808
rect 1454 5752 1459 5808
rect 0 5750 1459 5752
rect 0 5720 800 5750
rect 1393 5747 1459 5750
rect 2485 5472 2805 5473
rect 2485 5408 2493 5472
rect 2557 5408 2573 5472
rect 2637 5408 2653 5472
rect 2717 5408 2733 5472
rect 2797 5408 2805 5472
rect 2485 5407 2805 5408
rect 4027 5472 4347 5473
rect 4027 5408 4035 5472
rect 4099 5408 4115 5472
rect 4179 5408 4195 5472
rect 4259 5408 4275 5472
rect 4339 5408 4347 5472
rect 4027 5407 4347 5408
rect 5349 4994 5415 4997
rect 6033 4994 6833 5024
rect 5349 4992 6833 4994
rect 5349 4936 5354 4992
rect 5410 4936 6833 4992
rect 5349 4934 6833 4936
rect 5349 4931 5415 4934
rect 1715 4928 2035 4929
rect 1715 4864 1723 4928
rect 1787 4864 1803 4928
rect 1867 4864 1883 4928
rect 1947 4864 1963 4928
rect 2027 4864 2035 4928
rect 1715 4863 2035 4864
rect 3256 4928 3576 4929
rect 3256 4864 3264 4928
rect 3328 4864 3344 4928
rect 3408 4864 3424 4928
rect 3488 4864 3504 4928
rect 3568 4864 3576 4928
rect 3256 4863 3576 4864
rect 4798 4928 5118 4929
rect 4798 4864 4806 4928
rect 4870 4864 4886 4928
rect 4950 4864 4966 4928
rect 5030 4864 5046 4928
rect 5110 4864 5118 4928
rect 6033 4904 6833 4934
rect 4798 4863 5118 4864
rect 2485 4384 2805 4385
rect 2485 4320 2493 4384
rect 2557 4320 2573 4384
rect 2637 4320 2653 4384
rect 2717 4320 2733 4384
rect 2797 4320 2805 4384
rect 2485 4319 2805 4320
rect 4027 4384 4347 4385
rect 4027 4320 4035 4384
rect 4099 4320 4115 4384
rect 4179 4320 4195 4384
rect 4259 4320 4275 4384
rect 4339 4320 4347 4384
rect 4027 4319 4347 4320
rect 1715 3840 2035 3841
rect 1715 3776 1723 3840
rect 1787 3776 1803 3840
rect 1867 3776 1883 3840
rect 1947 3776 1963 3840
rect 2027 3776 2035 3840
rect 1715 3775 2035 3776
rect 3256 3840 3576 3841
rect 3256 3776 3264 3840
rect 3328 3776 3344 3840
rect 3408 3776 3424 3840
rect 3488 3776 3504 3840
rect 3568 3776 3576 3840
rect 3256 3775 3576 3776
rect 4798 3840 5118 3841
rect 4798 3776 4806 3840
rect 4870 3776 4886 3840
rect 4950 3776 4966 3840
rect 5030 3776 5046 3840
rect 5110 3776 5118 3840
rect 4798 3775 5118 3776
rect 2485 3296 2805 3297
rect 2485 3232 2493 3296
rect 2557 3232 2573 3296
rect 2637 3232 2653 3296
rect 2717 3232 2733 3296
rect 2797 3232 2805 3296
rect 2485 3231 2805 3232
rect 4027 3296 4347 3297
rect 4027 3232 4035 3296
rect 4099 3232 4115 3296
rect 4179 3232 4195 3296
rect 4259 3232 4275 3296
rect 4339 3232 4347 3296
rect 4027 3231 4347 3232
rect 0 2818 800 2848
rect 1393 2818 1459 2821
rect 0 2816 1459 2818
rect 0 2760 1398 2816
rect 1454 2760 1459 2816
rect 0 2758 1459 2760
rect 0 2728 800 2758
rect 1393 2755 1459 2758
rect 1715 2752 2035 2753
rect 1715 2688 1723 2752
rect 1787 2688 1803 2752
rect 1867 2688 1883 2752
rect 1947 2688 1963 2752
rect 2027 2688 2035 2752
rect 1715 2687 2035 2688
rect 3256 2752 3576 2753
rect 3256 2688 3264 2752
rect 3328 2688 3344 2752
rect 3408 2688 3424 2752
rect 3488 2688 3504 2752
rect 3568 2688 3576 2752
rect 3256 2687 3576 2688
rect 4798 2752 5118 2753
rect 4798 2688 4806 2752
rect 4870 2688 4886 2752
rect 4950 2688 4966 2752
rect 5030 2688 5046 2752
rect 5110 2688 5118 2752
rect 4798 2687 5118 2688
rect 4061 2410 4127 2413
rect 4061 2408 5090 2410
rect 4061 2352 4066 2408
rect 4122 2352 5090 2408
rect 4061 2350 5090 2352
rect 4061 2347 4127 2350
rect 2485 2208 2805 2209
rect 2485 2144 2493 2208
rect 2557 2144 2573 2208
rect 2637 2144 2653 2208
rect 2717 2144 2733 2208
rect 2797 2144 2805 2208
rect 2485 2143 2805 2144
rect 4027 2208 4347 2209
rect 4027 2144 4035 2208
rect 4099 2144 4115 2208
rect 4179 2144 4195 2208
rect 4259 2144 4275 2208
rect 4339 2144 4347 2208
rect 4027 2143 4347 2144
rect 5030 2002 5090 2350
rect 6033 2002 6833 2032
rect 5030 1942 6833 2002
rect 6033 1912 6833 1942
<< via3 >>
rect 2493 8732 2557 8736
rect 2493 8676 2497 8732
rect 2497 8676 2553 8732
rect 2553 8676 2557 8732
rect 2493 8672 2557 8676
rect 2573 8732 2637 8736
rect 2573 8676 2577 8732
rect 2577 8676 2633 8732
rect 2633 8676 2637 8732
rect 2573 8672 2637 8676
rect 2653 8732 2717 8736
rect 2653 8676 2657 8732
rect 2657 8676 2713 8732
rect 2713 8676 2717 8732
rect 2653 8672 2717 8676
rect 2733 8732 2797 8736
rect 2733 8676 2737 8732
rect 2737 8676 2793 8732
rect 2793 8676 2797 8732
rect 2733 8672 2797 8676
rect 4035 8732 4099 8736
rect 4035 8676 4039 8732
rect 4039 8676 4095 8732
rect 4095 8676 4099 8732
rect 4035 8672 4099 8676
rect 4115 8732 4179 8736
rect 4115 8676 4119 8732
rect 4119 8676 4175 8732
rect 4175 8676 4179 8732
rect 4115 8672 4179 8676
rect 4195 8732 4259 8736
rect 4195 8676 4199 8732
rect 4199 8676 4255 8732
rect 4255 8676 4259 8732
rect 4195 8672 4259 8676
rect 4275 8732 4339 8736
rect 4275 8676 4279 8732
rect 4279 8676 4335 8732
rect 4335 8676 4339 8732
rect 4275 8672 4339 8676
rect 1723 8188 1787 8192
rect 1723 8132 1727 8188
rect 1727 8132 1783 8188
rect 1783 8132 1787 8188
rect 1723 8128 1787 8132
rect 1803 8188 1867 8192
rect 1803 8132 1807 8188
rect 1807 8132 1863 8188
rect 1863 8132 1867 8188
rect 1803 8128 1867 8132
rect 1883 8188 1947 8192
rect 1883 8132 1887 8188
rect 1887 8132 1943 8188
rect 1943 8132 1947 8188
rect 1883 8128 1947 8132
rect 1963 8188 2027 8192
rect 1963 8132 1967 8188
rect 1967 8132 2023 8188
rect 2023 8132 2027 8188
rect 1963 8128 2027 8132
rect 3264 8188 3328 8192
rect 3264 8132 3268 8188
rect 3268 8132 3324 8188
rect 3324 8132 3328 8188
rect 3264 8128 3328 8132
rect 3344 8188 3408 8192
rect 3344 8132 3348 8188
rect 3348 8132 3404 8188
rect 3404 8132 3408 8188
rect 3344 8128 3408 8132
rect 3424 8188 3488 8192
rect 3424 8132 3428 8188
rect 3428 8132 3484 8188
rect 3484 8132 3488 8188
rect 3424 8128 3488 8132
rect 3504 8188 3568 8192
rect 3504 8132 3508 8188
rect 3508 8132 3564 8188
rect 3564 8132 3568 8188
rect 3504 8128 3568 8132
rect 4806 8188 4870 8192
rect 4806 8132 4810 8188
rect 4810 8132 4866 8188
rect 4866 8132 4870 8188
rect 4806 8128 4870 8132
rect 4886 8188 4950 8192
rect 4886 8132 4890 8188
rect 4890 8132 4946 8188
rect 4946 8132 4950 8188
rect 4886 8128 4950 8132
rect 4966 8188 5030 8192
rect 4966 8132 4970 8188
rect 4970 8132 5026 8188
rect 5026 8132 5030 8188
rect 4966 8128 5030 8132
rect 5046 8188 5110 8192
rect 5046 8132 5050 8188
rect 5050 8132 5106 8188
rect 5106 8132 5110 8188
rect 5046 8128 5110 8132
rect 2493 7644 2557 7648
rect 2493 7588 2497 7644
rect 2497 7588 2553 7644
rect 2553 7588 2557 7644
rect 2493 7584 2557 7588
rect 2573 7644 2637 7648
rect 2573 7588 2577 7644
rect 2577 7588 2633 7644
rect 2633 7588 2637 7644
rect 2573 7584 2637 7588
rect 2653 7644 2717 7648
rect 2653 7588 2657 7644
rect 2657 7588 2713 7644
rect 2713 7588 2717 7644
rect 2653 7584 2717 7588
rect 2733 7644 2797 7648
rect 2733 7588 2737 7644
rect 2737 7588 2793 7644
rect 2793 7588 2797 7644
rect 2733 7584 2797 7588
rect 4035 7644 4099 7648
rect 4035 7588 4039 7644
rect 4039 7588 4095 7644
rect 4095 7588 4099 7644
rect 4035 7584 4099 7588
rect 4115 7644 4179 7648
rect 4115 7588 4119 7644
rect 4119 7588 4175 7644
rect 4175 7588 4179 7644
rect 4115 7584 4179 7588
rect 4195 7644 4259 7648
rect 4195 7588 4199 7644
rect 4199 7588 4255 7644
rect 4255 7588 4259 7644
rect 4195 7584 4259 7588
rect 4275 7644 4339 7648
rect 4275 7588 4279 7644
rect 4279 7588 4335 7644
rect 4335 7588 4339 7644
rect 4275 7584 4339 7588
rect 1723 7100 1787 7104
rect 1723 7044 1727 7100
rect 1727 7044 1783 7100
rect 1783 7044 1787 7100
rect 1723 7040 1787 7044
rect 1803 7100 1867 7104
rect 1803 7044 1807 7100
rect 1807 7044 1863 7100
rect 1863 7044 1867 7100
rect 1803 7040 1867 7044
rect 1883 7100 1947 7104
rect 1883 7044 1887 7100
rect 1887 7044 1943 7100
rect 1943 7044 1947 7100
rect 1883 7040 1947 7044
rect 1963 7100 2027 7104
rect 1963 7044 1967 7100
rect 1967 7044 2023 7100
rect 2023 7044 2027 7100
rect 1963 7040 2027 7044
rect 3264 7100 3328 7104
rect 3264 7044 3268 7100
rect 3268 7044 3324 7100
rect 3324 7044 3328 7100
rect 3264 7040 3328 7044
rect 3344 7100 3408 7104
rect 3344 7044 3348 7100
rect 3348 7044 3404 7100
rect 3404 7044 3408 7100
rect 3344 7040 3408 7044
rect 3424 7100 3488 7104
rect 3424 7044 3428 7100
rect 3428 7044 3484 7100
rect 3484 7044 3488 7100
rect 3424 7040 3488 7044
rect 3504 7100 3568 7104
rect 3504 7044 3508 7100
rect 3508 7044 3564 7100
rect 3564 7044 3568 7100
rect 3504 7040 3568 7044
rect 4806 7100 4870 7104
rect 4806 7044 4810 7100
rect 4810 7044 4866 7100
rect 4866 7044 4870 7100
rect 4806 7040 4870 7044
rect 4886 7100 4950 7104
rect 4886 7044 4890 7100
rect 4890 7044 4946 7100
rect 4946 7044 4950 7100
rect 4886 7040 4950 7044
rect 4966 7100 5030 7104
rect 4966 7044 4970 7100
rect 4970 7044 5026 7100
rect 5026 7044 5030 7100
rect 4966 7040 5030 7044
rect 5046 7100 5110 7104
rect 5046 7044 5050 7100
rect 5050 7044 5106 7100
rect 5106 7044 5110 7100
rect 5046 7040 5110 7044
rect 2493 6556 2557 6560
rect 2493 6500 2497 6556
rect 2497 6500 2553 6556
rect 2553 6500 2557 6556
rect 2493 6496 2557 6500
rect 2573 6556 2637 6560
rect 2573 6500 2577 6556
rect 2577 6500 2633 6556
rect 2633 6500 2637 6556
rect 2573 6496 2637 6500
rect 2653 6556 2717 6560
rect 2653 6500 2657 6556
rect 2657 6500 2713 6556
rect 2713 6500 2717 6556
rect 2653 6496 2717 6500
rect 2733 6556 2797 6560
rect 2733 6500 2737 6556
rect 2737 6500 2793 6556
rect 2793 6500 2797 6556
rect 2733 6496 2797 6500
rect 4035 6556 4099 6560
rect 4035 6500 4039 6556
rect 4039 6500 4095 6556
rect 4095 6500 4099 6556
rect 4035 6496 4099 6500
rect 4115 6556 4179 6560
rect 4115 6500 4119 6556
rect 4119 6500 4175 6556
rect 4175 6500 4179 6556
rect 4115 6496 4179 6500
rect 4195 6556 4259 6560
rect 4195 6500 4199 6556
rect 4199 6500 4255 6556
rect 4255 6500 4259 6556
rect 4195 6496 4259 6500
rect 4275 6556 4339 6560
rect 4275 6500 4279 6556
rect 4279 6500 4335 6556
rect 4335 6500 4339 6556
rect 4275 6496 4339 6500
rect 1723 6012 1787 6016
rect 1723 5956 1727 6012
rect 1727 5956 1783 6012
rect 1783 5956 1787 6012
rect 1723 5952 1787 5956
rect 1803 6012 1867 6016
rect 1803 5956 1807 6012
rect 1807 5956 1863 6012
rect 1863 5956 1867 6012
rect 1803 5952 1867 5956
rect 1883 6012 1947 6016
rect 1883 5956 1887 6012
rect 1887 5956 1943 6012
rect 1943 5956 1947 6012
rect 1883 5952 1947 5956
rect 1963 6012 2027 6016
rect 1963 5956 1967 6012
rect 1967 5956 2023 6012
rect 2023 5956 2027 6012
rect 1963 5952 2027 5956
rect 3264 6012 3328 6016
rect 3264 5956 3268 6012
rect 3268 5956 3324 6012
rect 3324 5956 3328 6012
rect 3264 5952 3328 5956
rect 3344 6012 3408 6016
rect 3344 5956 3348 6012
rect 3348 5956 3404 6012
rect 3404 5956 3408 6012
rect 3344 5952 3408 5956
rect 3424 6012 3488 6016
rect 3424 5956 3428 6012
rect 3428 5956 3484 6012
rect 3484 5956 3488 6012
rect 3424 5952 3488 5956
rect 3504 6012 3568 6016
rect 3504 5956 3508 6012
rect 3508 5956 3564 6012
rect 3564 5956 3568 6012
rect 3504 5952 3568 5956
rect 4806 6012 4870 6016
rect 4806 5956 4810 6012
rect 4810 5956 4866 6012
rect 4866 5956 4870 6012
rect 4806 5952 4870 5956
rect 4886 6012 4950 6016
rect 4886 5956 4890 6012
rect 4890 5956 4946 6012
rect 4946 5956 4950 6012
rect 4886 5952 4950 5956
rect 4966 6012 5030 6016
rect 4966 5956 4970 6012
rect 4970 5956 5026 6012
rect 5026 5956 5030 6012
rect 4966 5952 5030 5956
rect 5046 6012 5110 6016
rect 5046 5956 5050 6012
rect 5050 5956 5106 6012
rect 5106 5956 5110 6012
rect 5046 5952 5110 5956
rect 2493 5468 2557 5472
rect 2493 5412 2497 5468
rect 2497 5412 2553 5468
rect 2553 5412 2557 5468
rect 2493 5408 2557 5412
rect 2573 5468 2637 5472
rect 2573 5412 2577 5468
rect 2577 5412 2633 5468
rect 2633 5412 2637 5468
rect 2573 5408 2637 5412
rect 2653 5468 2717 5472
rect 2653 5412 2657 5468
rect 2657 5412 2713 5468
rect 2713 5412 2717 5468
rect 2653 5408 2717 5412
rect 2733 5468 2797 5472
rect 2733 5412 2737 5468
rect 2737 5412 2793 5468
rect 2793 5412 2797 5468
rect 2733 5408 2797 5412
rect 4035 5468 4099 5472
rect 4035 5412 4039 5468
rect 4039 5412 4095 5468
rect 4095 5412 4099 5468
rect 4035 5408 4099 5412
rect 4115 5468 4179 5472
rect 4115 5412 4119 5468
rect 4119 5412 4175 5468
rect 4175 5412 4179 5468
rect 4115 5408 4179 5412
rect 4195 5468 4259 5472
rect 4195 5412 4199 5468
rect 4199 5412 4255 5468
rect 4255 5412 4259 5468
rect 4195 5408 4259 5412
rect 4275 5468 4339 5472
rect 4275 5412 4279 5468
rect 4279 5412 4335 5468
rect 4335 5412 4339 5468
rect 4275 5408 4339 5412
rect 1723 4924 1787 4928
rect 1723 4868 1727 4924
rect 1727 4868 1783 4924
rect 1783 4868 1787 4924
rect 1723 4864 1787 4868
rect 1803 4924 1867 4928
rect 1803 4868 1807 4924
rect 1807 4868 1863 4924
rect 1863 4868 1867 4924
rect 1803 4864 1867 4868
rect 1883 4924 1947 4928
rect 1883 4868 1887 4924
rect 1887 4868 1943 4924
rect 1943 4868 1947 4924
rect 1883 4864 1947 4868
rect 1963 4924 2027 4928
rect 1963 4868 1967 4924
rect 1967 4868 2023 4924
rect 2023 4868 2027 4924
rect 1963 4864 2027 4868
rect 3264 4924 3328 4928
rect 3264 4868 3268 4924
rect 3268 4868 3324 4924
rect 3324 4868 3328 4924
rect 3264 4864 3328 4868
rect 3344 4924 3408 4928
rect 3344 4868 3348 4924
rect 3348 4868 3404 4924
rect 3404 4868 3408 4924
rect 3344 4864 3408 4868
rect 3424 4924 3488 4928
rect 3424 4868 3428 4924
rect 3428 4868 3484 4924
rect 3484 4868 3488 4924
rect 3424 4864 3488 4868
rect 3504 4924 3568 4928
rect 3504 4868 3508 4924
rect 3508 4868 3564 4924
rect 3564 4868 3568 4924
rect 3504 4864 3568 4868
rect 4806 4924 4870 4928
rect 4806 4868 4810 4924
rect 4810 4868 4866 4924
rect 4866 4868 4870 4924
rect 4806 4864 4870 4868
rect 4886 4924 4950 4928
rect 4886 4868 4890 4924
rect 4890 4868 4946 4924
rect 4946 4868 4950 4924
rect 4886 4864 4950 4868
rect 4966 4924 5030 4928
rect 4966 4868 4970 4924
rect 4970 4868 5026 4924
rect 5026 4868 5030 4924
rect 4966 4864 5030 4868
rect 5046 4924 5110 4928
rect 5046 4868 5050 4924
rect 5050 4868 5106 4924
rect 5106 4868 5110 4924
rect 5046 4864 5110 4868
rect 2493 4380 2557 4384
rect 2493 4324 2497 4380
rect 2497 4324 2553 4380
rect 2553 4324 2557 4380
rect 2493 4320 2557 4324
rect 2573 4380 2637 4384
rect 2573 4324 2577 4380
rect 2577 4324 2633 4380
rect 2633 4324 2637 4380
rect 2573 4320 2637 4324
rect 2653 4380 2717 4384
rect 2653 4324 2657 4380
rect 2657 4324 2713 4380
rect 2713 4324 2717 4380
rect 2653 4320 2717 4324
rect 2733 4380 2797 4384
rect 2733 4324 2737 4380
rect 2737 4324 2793 4380
rect 2793 4324 2797 4380
rect 2733 4320 2797 4324
rect 4035 4380 4099 4384
rect 4035 4324 4039 4380
rect 4039 4324 4095 4380
rect 4095 4324 4099 4380
rect 4035 4320 4099 4324
rect 4115 4380 4179 4384
rect 4115 4324 4119 4380
rect 4119 4324 4175 4380
rect 4175 4324 4179 4380
rect 4115 4320 4179 4324
rect 4195 4380 4259 4384
rect 4195 4324 4199 4380
rect 4199 4324 4255 4380
rect 4255 4324 4259 4380
rect 4195 4320 4259 4324
rect 4275 4380 4339 4384
rect 4275 4324 4279 4380
rect 4279 4324 4335 4380
rect 4335 4324 4339 4380
rect 4275 4320 4339 4324
rect 1723 3836 1787 3840
rect 1723 3780 1727 3836
rect 1727 3780 1783 3836
rect 1783 3780 1787 3836
rect 1723 3776 1787 3780
rect 1803 3836 1867 3840
rect 1803 3780 1807 3836
rect 1807 3780 1863 3836
rect 1863 3780 1867 3836
rect 1803 3776 1867 3780
rect 1883 3836 1947 3840
rect 1883 3780 1887 3836
rect 1887 3780 1943 3836
rect 1943 3780 1947 3836
rect 1883 3776 1947 3780
rect 1963 3836 2027 3840
rect 1963 3780 1967 3836
rect 1967 3780 2023 3836
rect 2023 3780 2027 3836
rect 1963 3776 2027 3780
rect 3264 3836 3328 3840
rect 3264 3780 3268 3836
rect 3268 3780 3324 3836
rect 3324 3780 3328 3836
rect 3264 3776 3328 3780
rect 3344 3836 3408 3840
rect 3344 3780 3348 3836
rect 3348 3780 3404 3836
rect 3404 3780 3408 3836
rect 3344 3776 3408 3780
rect 3424 3836 3488 3840
rect 3424 3780 3428 3836
rect 3428 3780 3484 3836
rect 3484 3780 3488 3836
rect 3424 3776 3488 3780
rect 3504 3836 3568 3840
rect 3504 3780 3508 3836
rect 3508 3780 3564 3836
rect 3564 3780 3568 3836
rect 3504 3776 3568 3780
rect 4806 3836 4870 3840
rect 4806 3780 4810 3836
rect 4810 3780 4866 3836
rect 4866 3780 4870 3836
rect 4806 3776 4870 3780
rect 4886 3836 4950 3840
rect 4886 3780 4890 3836
rect 4890 3780 4946 3836
rect 4946 3780 4950 3836
rect 4886 3776 4950 3780
rect 4966 3836 5030 3840
rect 4966 3780 4970 3836
rect 4970 3780 5026 3836
rect 5026 3780 5030 3836
rect 4966 3776 5030 3780
rect 5046 3836 5110 3840
rect 5046 3780 5050 3836
rect 5050 3780 5106 3836
rect 5106 3780 5110 3836
rect 5046 3776 5110 3780
rect 2493 3292 2557 3296
rect 2493 3236 2497 3292
rect 2497 3236 2553 3292
rect 2553 3236 2557 3292
rect 2493 3232 2557 3236
rect 2573 3292 2637 3296
rect 2573 3236 2577 3292
rect 2577 3236 2633 3292
rect 2633 3236 2637 3292
rect 2573 3232 2637 3236
rect 2653 3292 2717 3296
rect 2653 3236 2657 3292
rect 2657 3236 2713 3292
rect 2713 3236 2717 3292
rect 2653 3232 2717 3236
rect 2733 3292 2797 3296
rect 2733 3236 2737 3292
rect 2737 3236 2793 3292
rect 2793 3236 2797 3292
rect 2733 3232 2797 3236
rect 4035 3292 4099 3296
rect 4035 3236 4039 3292
rect 4039 3236 4095 3292
rect 4095 3236 4099 3292
rect 4035 3232 4099 3236
rect 4115 3292 4179 3296
rect 4115 3236 4119 3292
rect 4119 3236 4175 3292
rect 4175 3236 4179 3292
rect 4115 3232 4179 3236
rect 4195 3292 4259 3296
rect 4195 3236 4199 3292
rect 4199 3236 4255 3292
rect 4255 3236 4259 3292
rect 4195 3232 4259 3236
rect 4275 3292 4339 3296
rect 4275 3236 4279 3292
rect 4279 3236 4335 3292
rect 4335 3236 4339 3292
rect 4275 3232 4339 3236
rect 1723 2748 1787 2752
rect 1723 2692 1727 2748
rect 1727 2692 1783 2748
rect 1783 2692 1787 2748
rect 1723 2688 1787 2692
rect 1803 2748 1867 2752
rect 1803 2692 1807 2748
rect 1807 2692 1863 2748
rect 1863 2692 1867 2748
rect 1803 2688 1867 2692
rect 1883 2748 1947 2752
rect 1883 2692 1887 2748
rect 1887 2692 1943 2748
rect 1943 2692 1947 2748
rect 1883 2688 1947 2692
rect 1963 2748 2027 2752
rect 1963 2692 1967 2748
rect 1967 2692 2023 2748
rect 2023 2692 2027 2748
rect 1963 2688 2027 2692
rect 3264 2748 3328 2752
rect 3264 2692 3268 2748
rect 3268 2692 3324 2748
rect 3324 2692 3328 2748
rect 3264 2688 3328 2692
rect 3344 2748 3408 2752
rect 3344 2692 3348 2748
rect 3348 2692 3404 2748
rect 3404 2692 3408 2748
rect 3344 2688 3408 2692
rect 3424 2748 3488 2752
rect 3424 2692 3428 2748
rect 3428 2692 3484 2748
rect 3484 2692 3488 2748
rect 3424 2688 3488 2692
rect 3504 2748 3568 2752
rect 3504 2692 3508 2748
rect 3508 2692 3564 2748
rect 3564 2692 3568 2748
rect 3504 2688 3568 2692
rect 4806 2748 4870 2752
rect 4806 2692 4810 2748
rect 4810 2692 4866 2748
rect 4866 2692 4870 2748
rect 4806 2688 4870 2692
rect 4886 2748 4950 2752
rect 4886 2692 4890 2748
rect 4890 2692 4946 2748
rect 4946 2692 4950 2748
rect 4886 2688 4950 2692
rect 4966 2748 5030 2752
rect 4966 2692 4970 2748
rect 4970 2692 5026 2748
rect 5026 2692 5030 2748
rect 4966 2688 5030 2692
rect 5046 2748 5110 2752
rect 5046 2692 5050 2748
rect 5050 2692 5106 2748
rect 5106 2692 5110 2748
rect 5046 2688 5110 2692
rect 2493 2204 2557 2208
rect 2493 2148 2497 2204
rect 2497 2148 2553 2204
rect 2553 2148 2557 2204
rect 2493 2144 2557 2148
rect 2573 2204 2637 2208
rect 2573 2148 2577 2204
rect 2577 2148 2633 2204
rect 2633 2148 2637 2204
rect 2573 2144 2637 2148
rect 2653 2204 2717 2208
rect 2653 2148 2657 2204
rect 2657 2148 2713 2204
rect 2713 2148 2717 2204
rect 2653 2144 2717 2148
rect 2733 2204 2797 2208
rect 2733 2148 2737 2204
rect 2737 2148 2793 2204
rect 2793 2148 2797 2204
rect 2733 2144 2797 2148
rect 4035 2204 4099 2208
rect 4035 2148 4039 2204
rect 4039 2148 4095 2204
rect 4095 2148 4099 2204
rect 4035 2144 4099 2148
rect 4115 2204 4179 2208
rect 4115 2148 4119 2204
rect 4119 2148 4175 2204
rect 4175 2148 4179 2204
rect 4115 2144 4179 2148
rect 4195 2204 4259 2208
rect 4195 2148 4199 2204
rect 4199 2148 4255 2204
rect 4255 2148 4259 2204
rect 4195 2144 4259 2148
rect 4275 2204 4339 2208
rect 4275 2148 4279 2204
rect 4279 2148 4335 2204
rect 4335 2148 4339 2204
rect 4275 2144 4339 2148
<< metal4 >>
rect 1715 8192 2035 8752
rect 1715 8128 1723 8192
rect 1787 8128 1803 8192
rect 1867 8128 1883 8192
rect 1947 8128 1963 8192
rect 2027 8128 2035 8192
rect 1715 7767 2035 8128
rect 1715 7531 1757 7767
rect 1993 7531 2035 7767
rect 1715 7104 2035 7531
rect 1715 7040 1723 7104
rect 1787 7040 1803 7104
rect 1867 7040 1883 7104
rect 1947 7040 1963 7104
rect 2027 7040 2035 7104
rect 1715 6016 2035 7040
rect 1715 5952 1723 6016
rect 1787 5952 1803 6016
rect 1867 5952 1883 6016
rect 1947 5952 1963 6016
rect 2027 5952 2035 6016
rect 1715 5558 2035 5952
rect 1715 5322 1757 5558
rect 1993 5322 2035 5558
rect 1715 4928 2035 5322
rect 1715 4864 1723 4928
rect 1787 4864 1803 4928
rect 1867 4864 1883 4928
rect 1947 4864 1963 4928
rect 2027 4864 2035 4928
rect 1715 3840 2035 4864
rect 1715 3776 1723 3840
rect 1787 3776 1803 3840
rect 1867 3776 1883 3840
rect 1947 3776 1963 3840
rect 2027 3776 2035 3840
rect 1715 3350 2035 3776
rect 1715 3114 1757 3350
rect 1993 3114 2035 3350
rect 1715 2752 2035 3114
rect 1715 2688 1723 2752
rect 1787 2688 1803 2752
rect 1867 2688 1883 2752
rect 1947 2688 1963 2752
rect 2027 2688 2035 2752
rect 1715 2128 2035 2688
rect 2485 8736 2805 8752
rect 2485 8672 2493 8736
rect 2557 8672 2573 8736
rect 2637 8672 2653 8736
rect 2717 8672 2733 8736
rect 2797 8672 2805 8736
rect 2485 7648 2805 8672
rect 2485 7584 2493 7648
rect 2557 7584 2573 7648
rect 2637 7584 2653 7648
rect 2717 7584 2733 7648
rect 2797 7584 2805 7648
rect 2485 6663 2805 7584
rect 2485 6560 2527 6663
rect 2763 6560 2805 6663
rect 2485 6496 2493 6560
rect 2797 6496 2805 6560
rect 2485 6427 2527 6496
rect 2763 6427 2805 6496
rect 2485 5472 2805 6427
rect 2485 5408 2493 5472
rect 2557 5408 2573 5472
rect 2637 5408 2653 5472
rect 2717 5408 2733 5472
rect 2797 5408 2805 5472
rect 2485 4454 2805 5408
rect 2485 4384 2527 4454
rect 2763 4384 2805 4454
rect 2485 4320 2493 4384
rect 2797 4320 2805 4384
rect 2485 4218 2527 4320
rect 2763 4218 2805 4320
rect 2485 3296 2805 4218
rect 2485 3232 2493 3296
rect 2557 3232 2573 3296
rect 2637 3232 2653 3296
rect 2717 3232 2733 3296
rect 2797 3232 2805 3296
rect 2485 2208 2805 3232
rect 2485 2144 2493 2208
rect 2557 2144 2573 2208
rect 2637 2144 2653 2208
rect 2717 2144 2733 2208
rect 2797 2144 2805 2208
rect 2485 2128 2805 2144
rect 3256 8192 3576 8752
rect 3256 8128 3264 8192
rect 3328 8128 3344 8192
rect 3408 8128 3424 8192
rect 3488 8128 3504 8192
rect 3568 8128 3576 8192
rect 3256 7767 3576 8128
rect 3256 7531 3298 7767
rect 3534 7531 3576 7767
rect 3256 7104 3576 7531
rect 3256 7040 3264 7104
rect 3328 7040 3344 7104
rect 3408 7040 3424 7104
rect 3488 7040 3504 7104
rect 3568 7040 3576 7104
rect 3256 6016 3576 7040
rect 3256 5952 3264 6016
rect 3328 5952 3344 6016
rect 3408 5952 3424 6016
rect 3488 5952 3504 6016
rect 3568 5952 3576 6016
rect 3256 5558 3576 5952
rect 3256 5322 3298 5558
rect 3534 5322 3576 5558
rect 3256 4928 3576 5322
rect 3256 4864 3264 4928
rect 3328 4864 3344 4928
rect 3408 4864 3424 4928
rect 3488 4864 3504 4928
rect 3568 4864 3576 4928
rect 3256 3840 3576 4864
rect 3256 3776 3264 3840
rect 3328 3776 3344 3840
rect 3408 3776 3424 3840
rect 3488 3776 3504 3840
rect 3568 3776 3576 3840
rect 3256 3350 3576 3776
rect 3256 3114 3298 3350
rect 3534 3114 3576 3350
rect 3256 2752 3576 3114
rect 3256 2688 3264 2752
rect 3328 2688 3344 2752
rect 3408 2688 3424 2752
rect 3488 2688 3504 2752
rect 3568 2688 3576 2752
rect 3256 2128 3576 2688
rect 4027 8736 4347 8752
rect 4027 8672 4035 8736
rect 4099 8672 4115 8736
rect 4179 8672 4195 8736
rect 4259 8672 4275 8736
rect 4339 8672 4347 8736
rect 4027 7648 4347 8672
rect 4027 7584 4035 7648
rect 4099 7584 4115 7648
rect 4179 7584 4195 7648
rect 4259 7584 4275 7648
rect 4339 7584 4347 7648
rect 4027 6663 4347 7584
rect 4027 6560 4069 6663
rect 4305 6560 4347 6663
rect 4027 6496 4035 6560
rect 4339 6496 4347 6560
rect 4027 6427 4069 6496
rect 4305 6427 4347 6496
rect 4027 5472 4347 6427
rect 4027 5408 4035 5472
rect 4099 5408 4115 5472
rect 4179 5408 4195 5472
rect 4259 5408 4275 5472
rect 4339 5408 4347 5472
rect 4027 4454 4347 5408
rect 4027 4384 4069 4454
rect 4305 4384 4347 4454
rect 4027 4320 4035 4384
rect 4339 4320 4347 4384
rect 4027 4218 4069 4320
rect 4305 4218 4347 4320
rect 4027 3296 4347 4218
rect 4027 3232 4035 3296
rect 4099 3232 4115 3296
rect 4179 3232 4195 3296
rect 4259 3232 4275 3296
rect 4339 3232 4347 3296
rect 4027 2208 4347 3232
rect 4027 2144 4035 2208
rect 4099 2144 4115 2208
rect 4179 2144 4195 2208
rect 4259 2144 4275 2208
rect 4339 2144 4347 2208
rect 4027 2128 4347 2144
rect 4798 8192 5118 8752
rect 4798 8128 4806 8192
rect 4870 8128 4886 8192
rect 4950 8128 4966 8192
rect 5030 8128 5046 8192
rect 5110 8128 5118 8192
rect 4798 7767 5118 8128
rect 4798 7531 4840 7767
rect 5076 7531 5118 7767
rect 4798 7104 5118 7531
rect 4798 7040 4806 7104
rect 4870 7040 4886 7104
rect 4950 7040 4966 7104
rect 5030 7040 5046 7104
rect 5110 7040 5118 7104
rect 4798 6016 5118 7040
rect 4798 5952 4806 6016
rect 4870 5952 4886 6016
rect 4950 5952 4966 6016
rect 5030 5952 5046 6016
rect 5110 5952 5118 6016
rect 4798 5558 5118 5952
rect 4798 5322 4840 5558
rect 5076 5322 5118 5558
rect 4798 4928 5118 5322
rect 4798 4864 4806 4928
rect 4870 4864 4886 4928
rect 4950 4864 4966 4928
rect 5030 4864 5046 4928
rect 5110 4864 5118 4928
rect 4798 3840 5118 4864
rect 4798 3776 4806 3840
rect 4870 3776 4886 3840
rect 4950 3776 4966 3840
rect 5030 3776 5046 3840
rect 5110 3776 5118 3840
rect 4798 3350 5118 3776
rect 4798 3114 4840 3350
rect 5076 3114 5118 3350
rect 4798 2752 5118 3114
rect 4798 2688 4806 2752
rect 4870 2688 4886 2752
rect 4950 2688 4966 2752
rect 5030 2688 5046 2752
rect 5110 2688 5118 2752
rect 4798 2128 5118 2688
<< via4 >>
rect 1757 7531 1993 7767
rect 1757 5322 1993 5558
rect 1757 3114 1993 3350
rect 2527 6560 2763 6663
rect 2527 6496 2557 6560
rect 2557 6496 2573 6560
rect 2573 6496 2637 6560
rect 2637 6496 2653 6560
rect 2653 6496 2717 6560
rect 2717 6496 2733 6560
rect 2733 6496 2763 6560
rect 2527 6427 2763 6496
rect 2527 4384 2763 4454
rect 2527 4320 2557 4384
rect 2557 4320 2573 4384
rect 2573 4320 2637 4384
rect 2637 4320 2653 4384
rect 2653 4320 2717 4384
rect 2717 4320 2733 4384
rect 2733 4320 2763 4384
rect 2527 4218 2763 4320
rect 3298 7531 3534 7767
rect 3298 5322 3534 5558
rect 3298 3114 3534 3350
rect 4069 6560 4305 6663
rect 4069 6496 4099 6560
rect 4099 6496 4115 6560
rect 4115 6496 4179 6560
rect 4179 6496 4195 6560
rect 4195 6496 4259 6560
rect 4259 6496 4275 6560
rect 4275 6496 4305 6560
rect 4069 6427 4305 6496
rect 4069 4384 4305 4454
rect 4069 4320 4099 4384
rect 4099 4320 4115 4384
rect 4115 4320 4179 4384
rect 4179 4320 4195 4384
rect 4195 4320 4259 4384
rect 4259 4320 4275 4384
rect 4275 4320 4305 4384
rect 4069 4218 4305 4320
rect 4840 7531 5076 7767
rect 4840 5322 5076 5558
rect 4840 3114 5076 3350
<< metal5 >>
rect 1104 7767 5704 7809
rect 1104 7531 1757 7767
rect 1993 7531 3298 7767
rect 3534 7531 4840 7767
rect 5076 7531 5704 7767
rect 1104 7489 5704 7531
rect 1104 6663 5704 6705
rect 1104 6427 2527 6663
rect 2763 6427 4069 6663
rect 4305 6427 5704 6663
rect 1104 6385 5704 6427
rect 1104 5558 5704 5600
rect 1104 5322 1757 5558
rect 1993 5322 3298 5558
rect 3534 5322 4840 5558
rect 5076 5322 5704 5558
rect 1104 5280 5704 5322
rect 1104 4454 5704 4497
rect 1104 4218 2527 4454
rect 2763 4218 4069 4454
rect 4305 4218 5704 4454
rect 1104 4176 5704 4218
rect 1104 3350 5704 3392
rect 1104 3114 1757 3350
rect 1993 3114 3298 3350
rect 3534 3114 4840 3350
rect 5076 3114 5704 3350
rect 1104 3072 5704 3114
use sky130_fd_sc_hd__fill_1  FILLER_1_10 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1628835793
transform 1 0 2024 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_6 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1628835793
transform 1 0 1656 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1628835793
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1628835793
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _49_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1628835793
transform -1 0 2392 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input2 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1628835793
transform 1 0 1380 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input4 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1628835793
transform 1 0 1380 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13
timestamp 1628835793
transform 1 0 2300 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1628835793
transform 1 0 2944 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_1_14
timestamp 1628835793
transform 1 0 2392 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_21
timestamp 1628835793
transform 1 0 3036 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _52_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1628835793
transform 1 0 2760 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1628835793
transform -1 0 2944 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input7
timestamp 1628835793
transform -1 0 3680 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29
timestamp 1628835793
transform 1 0 3772 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_35
timestamp 1628835793
transform 1 0 4324 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_28
timestamp 1628835793
transform 1 0 3680 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_32
timestamp 1628835793
transform 1 0 4048 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_36
timestamp 1628835793
transform 1 0 4416 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_24 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1628835793
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp 1628835793
transform -1 0 4324 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input9
timestamp 1628835793
transform 1 0 4140 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_43
timestamp 1628835793
transform 1 0 5060 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_43
timestamp 1628835793
transform 1 0 5060 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1628835793
transform -1 0 5704 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1628835793
transform -1 0 5704 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _57_
timestamp 1628835793
transform 1 0 4784 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output11 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1628835793
transform 1 0 4692 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_3
timestamp 1628835793
transform 1 0 1380 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_7
timestamp 1628835793
transform 1 0 1748 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1628835793
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _44_
timestamp 1628835793
transform 1 0 1472 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__or3b_1  _53_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1628835793
transform -1 0 2760 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_2_18
timestamp 1628835793
transform 1 0 2760 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_26 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1628835793
transform 1 0 3496 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_2_32
timestamp 1628835793
transform 1 0 4048 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_25
timestamp 1628835793
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _41_
timestamp 1628835793
transform 1 0 3772 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_2_43
timestamp 1628835793
transform 1 0 5060 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1628835793
transform -1 0 5704 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input8
timestamp 1628835793
transform -1 0 5060 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_3
timestamp 1628835793
transform 1 0 1380 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_7
timestamp 1628835793
transform 1 0 1748 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1628835793
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__o41a_1  _54_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1628835793
transform 1 0 1840 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_3_17
timestamp 1628835793
transform 1 0 2668 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_25
timestamp 1628835793
transform 1 0 3404 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_29
timestamp 1628835793
transform 1 0 3772 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_33
timestamp 1628835793
transform 1 0 4140 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_37
timestamp 1628835793
transform 1 0 4508 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  _29_
timestamp 1628835793
transform 1 0 4232 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _37_
timestamp 1628835793
transform -1 0 3772 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_45
timestamp 1628835793
transform 1 0 5244 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1628835793
transform -1 0 5704 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_4_12
timestamp 1628835793
transform 1 0 2208 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1628835793
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__a2111o_1  _45_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1628835793
transform 1 0 1380 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_4_21 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1628835793
transform 1 0 3036 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _39_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1628835793
transform 1 0 2576 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp 1628835793
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_37
timestamp 1628835793
transform 1 0 4508 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_26
timestamp 1628835793
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__o2bb2a_1  _42_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1628835793
transform 1 0 3772 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_4_45
timestamp 1628835793
transform 1 0 5244 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1628835793
transform -1 0 5704 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_5_8
timestamp 1628835793
transform 1 0 1840 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1628835793
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _38_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1628835793
transform -1 0 1840 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__decap_8  FILLER_5_19
timestamp 1628835793
transform 1 0 2852 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _43_
timestamp 1628835793
transform -1 0 2852 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__decap_6  FILLER_5_32
timestamp 1628835793
transform 1 0 4048 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_38
timestamp 1628835793
transform 1 0 4600 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__or3_1  _36_
timestamp 1628835793
transform -1 0 4048 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__decap_4  FILLER_5_43
timestamp 1628835793
transform 1 0 5060 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1628835793
transform -1 0 5704 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output14
timestamp 1628835793
transform 1 0 4692 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_11
timestamp 1628835793
transform 1 0 2116 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_7
timestamp 1628835793
transform 1 0 1748 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_7_3
timestamp 1628835793
transform 1 0 1380 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1628835793
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1628835793
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _47_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1628835793
transform -1 0 1748 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__o22ai_1  _56_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1628835793
transform 1 0 1932 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__dlxtn_1  _60_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1628835793
transform 1 0 2208 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_24
timestamp 1628835793
transform 1 0 3312 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_14
timestamp 1628835793
transform 1 0 2392 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_22
timestamp 1628835793
transform 1 0 3128 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _40_
timestamp 1628835793
transform 1 0 2760 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_6_37
timestamp 1628835793
transform 1 0 4508 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_26
timestamp 1628835793
transform 1 0 3496 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_33
timestamp 1628835793
transform 1 0 4140 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_27
timestamp 1628835793
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _28_
timestamp 1628835793
transform 1 0 4508 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__a2bb2o_1  _35_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1628835793
transform 1 0 3772 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _46_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1628835793
transform -1 0 4140 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_6_45
timestamp 1628835793
transform 1 0 5244 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_7_40
timestamp 1628835793
transform 1 0 4784 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_46
timestamp 1628835793
transform 1 0 5336 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1628835793
transform -1 0 5704 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1628835793
transform -1 0 5704 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_8_6
timestamp 1628835793
transform 1 0 1656 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1628835793
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__o22ai_1  _55_
timestamp 1628835793
transform 1 0 2024 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  input3
timestamp 1628835793
transform 1 0 1380 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_8_15
timestamp 1628835793
transform 1 0 2484 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_23
timestamp 1628835793
transform 1 0 3220 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _48_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1628835793
transform -1 0 3220 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_27
timestamp 1628835793
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_34
timestamp 1628835793
transform 1 0 4232 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_38
timestamp 1628835793
transform 1 0 4600 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_28
timestamp 1628835793
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__or3_1  _34_
timestamp 1628835793
transform -1 0 4232 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__decap_4  FILLER_8_42
timestamp 1628835793
transform 1 0 4968 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_46
timestamp 1628835793
transform 1 0 5336 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1628835793
transform -1 0 5704 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input5
timestamp 1628835793
transform 1 0 4692 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_9_3
timestamp 1628835793
transform 1 0 1380 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1628835793
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__dlxtn_1  _59_
timestamp 1628835793
transform 1 0 1472 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_16
timestamp 1628835793
transform 1 0 2576 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__o41a_1  _51_
timestamp 1628835793
transform 1 0 2944 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_9_29
timestamp 1628835793
transform 1 0 3772 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__or4b_1  _50_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1628835793
transform -1 0 4876 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_9_41
timestamp 1628835793
transform 1 0 4876 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1628835793
transform -1 0 5704 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_10_3
timestamp 1628835793
transform 1 0 1380 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1628835793
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__dlxtn_1  _58_
timestamp 1628835793
transform -1 0 2852 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_19
timestamp 1628835793
transform 1 0 2852 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_27
timestamp 1628835793
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_36
timestamp 1628835793
transform 1 0 4416 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_29
timestamp 1628835793
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__o22a_1  _33_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1628835793
transform 1 0 3772 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_10_43
timestamp 1628835793
transform 1 0 5060 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1628835793
transform -1 0 5704 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _31_
timestamp 1628835793
transform -1 0 5060 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_11_7
timestamp 1628835793
transform 1 0 1748 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1628835793
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output12
timestamp 1628835793
transform -1 0 1748 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output13
timestamp 1628835793
transform -1 0 2484 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_11_15
timestamp 1628835793
transform 1 0 2484 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_11_24
timestamp 1628835793
transform 1 0 3312 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _32_
timestamp 1628835793
transform -1 0 3312 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_11_32
timestamp 1628835793
transform 1 0 4048 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_38
timestamp 1628835793
transform 1 0 4600 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_30
timestamp 1628835793
transform 1 0 3680 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _30_
timestamp 1628835793
transform -1 0 4048 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_11_43
timestamp 1628835793
transform 1 0 5060 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1628835793
transform -1 0 5704 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output10
timestamp 1628835793
transform 1 0 4692 0 -1 8704
box -38 -48 406 592
<< labels >>
rlabel metal5 s 1104 4177 5704 4497 6 VGND
port 0 nsew ground input
rlabel metal5 s 1104 3072 5704 3392 6 VPWR
port 1 nsew power input
rlabel metal2 s 2042 0 2098 800 6 en
port 2 nsew signal input
rlabel metal3 s 6033 7896 6833 8016 6 eno
port 3 nsew signal tristate
rlabel metal2 s 6090 0 6146 800 6 gs
port 4 nsew signal tristate
rlabel metal3 s 0 2728 800 2848 6 in[0]
port 5 nsew signal input
rlabel metal3 s 0 5720 800 5840 6 in[1]
port 6 nsew signal input
rlabel metal2 s 18 0 74 800 6 in[2]
port 7 nsew signal input
rlabel metal2 s 4618 10177 4674 10977 6 in[3]
port 8 nsew signal input
rlabel metal3 s 6033 1912 6833 2032 6 in[4]
port 9 nsew signal input
rlabel metal2 s 2594 10177 2650 10977 6 in[5]
port 10 nsew signal input
rlabel metal2 s 6642 10177 6698 10977 6 in[6]
port 11 nsew signal input
rlabel metal2 s 4066 0 4122 800 6 in[7]
port 12 nsew signal input
rlabel metal3 s 0 8712 800 8832 6 out[0]
port 13 nsew signal tristate
rlabel metal2 s 570 10177 626 10977 6 out[1]
port 14 nsew signal tristate
rlabel metal3 s 6033 4904 6833 5024 6 out[2]
port 15 nsew signal tristate
<< properties >>
string FIXED_BBOX 0 0 6833 10977
<< end >>
