magic
tech sky130A
magscale 1 2
timestamp 1629374143
<< obsli1 >>
rect 1104 2159 6043 8721
<< obsm1 >>
rect 14 2128 6702 8752
<< metal2 >>
rect 570 10177 626 10977
rect 2594 10177 2650 10977
rect 4618 10177 4674 10977
rect 6642 10177 6698 10977
rect 18 0 74 800
rect 2042 0 2098 800
rect 4066 0 4122 800
rect 6090 0 6146 800
<< obsm2 >>
rect 20 10121 514 10282
rect 682 10121 2538 10282
rect 2706 10121 4562 10282
rect 4730 10121 6586 10282
rect 20 856 6696 10121
rect 130 800 1986 856
rect 2154 800 4010 856
rect 4178 800 6034 856
rect 6202 800 6696 856
<< metal3 >>
rect 0 8712 800 8832
rect 6033 7896 6833 8016
rect 0 5720 800 5840
rect 6033 4904 6833 5024
rect 0 2728 800 2848
rect 6033 1912 6833 2032
<< obsm3 >>
rect 880 8632 6033 8805
rect 800 8096 6033 8632
rect 800 7816 5953 8096
rect 800 5920 6033 7816
rect 880 5640 6033 5920
rect 800 5104 6033 5640
rect 800 4824 5953 5104
rect 800 2928 6033 4824
rect 880 2648 6033 2928
rect 800 2112 6033 2648
rect 800 1942 5953 2112
<< obsm4 >>
rect 1715 2128 5118 8752
<< metal5 >>
rect 1104 4177 5704 4497
rect 1104 3072 5704 3392
<< obsm5 >>
rect 1104 4817 5704 7809
<< labels >>
rlabel metal5 s 1104 4177 5704 4497 6 VGND
port 1 nsew ground input
rlabel metal5 s 1104 3072 5704 3392 6 VPWR
port 2 nsew power input
rlabel metal2 s 2042 0 2098 800 6 en
port 3 nsew signal input
rlabel metal3 s 6033 7896 6833 8016 6 eno
port 4 nsew signal output
rlabel metal2 s 6090 0 6146 800 6 gs
port 5 nsew signal output
rlabel metal3 s 0 2728 800 2848 6 in[0]
port 6 nsew signal input
rlabel metal3 s 0 5720 800 5840 6 in[1]
port 7 nsew signal input
rlabel metal2 s 18 0 74 800 6 in[2]
port 8 nsew signal input
rlabel metal2 s 4618 10177 4674 10977 6 in[3]
port 9 nsew signal input
rlabel metal3 s 6033 1912 6833 2032 6 in[4]
port 10 nsew signal input
rlabel metal2 s 2594 10177 2650 10977 6 in[5]
port 11 nsew signal input
rlabel metal2 s 6642 10177 6698 10977 6 in[6]
port 12 nsew signal input
rlabel metal2 s 4066 0 4122 800 6 in[7]
port 13 nsew signal input
rlabel metal3 s 0 8712 800 8832 6 out[0]
port 14 nsew signal output
rlabel metal2 s 570 10177 626 10977 6 out[1]
port 15 nsew signal output
rlabel metal3 s 6033 4904 6833 5024 6 out[2]
port 16 nsew signal output
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 6833 10977
string LEFview TRUE
string GDS_FILE /openLANE_flow/designs/dvsd_pe/runs/run3/results/magic/dvsd_pe.gds
string GDS_END 268582
string GDS_START 135290
<< end >>

