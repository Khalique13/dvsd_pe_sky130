VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO dvsd_pe
  CLASS BLOCK ;
  FOREIGN dvsd_pe ;
  ORIGIN 0.000 0.000 ;
  SIZE 34.165 BY 54.885 ;
  PIN VGND
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 5.520 20.885 28.520 22.485 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 5.520 15.360 28.520 16.960 ;
    END
  END VPWR
  PIN en
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 10.210 0.000 10.490 4.000 ;
    END
  END en
  PIN eno
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 30.165 39.480 34.165 40.080 ;
    END
  END eno
  PIN gs
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 30.450 0.000 30.730 4.000 ;
    END
  END gs
  PIN in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 13.640 4.000 14.240 ;
    END
  END in[0]
  PIN in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 28.600 4.000 29.200 ;
    END
  END in[1]
  PIN in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.090 0.000 0.370 4.000 ;
    END
  END in[2]
  PIN in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 23.090 50.885 23.370 54.885 ;
    END
  END in[3]
  PIN in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 30.165 9.560 34.165 10.160 ;
    END
  END in[4]
  PIN in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.970 50.885 13.250 54.885 ;
    END
  END in[5]
  PIN in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 33.210 50.885 33.490 54.885 ;
    END
  END in[6]
  PIN in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 20.330 0.000 20.610 4.000 ;
    END
  END in[7]
  PIN out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 43.560 4.000 44.160 ;
    END
  END out[0]
  PIN out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2.850 50.885 3.130 54.885 ;
    END
  END out[1]
  PIN out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 30.165 24.520 34.165 25.120 ;
    END
  END out[2]
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 30.215 43.605 ;
      LAYER met1 ;
        RECT 0.070 10.640 33.510 43.760 ;
      LAYER met2 ;
        RECT 0.100 50.605 2.570 51.410 ;
        RECT 3.410 50.605 12.690 51.410 ;
        RECT 13.530 50.605 22.810 51.410 ;
        RECT 23.650 50.605 32.930 51.410 ;
        RECT 0.100 4.280 33.480 50.605 ;
        RECT 0.650 4.000 9.930 4.280 ;
        RECT 10.770 4.000 20.050 4.280 ;
        RECT 20.890 4.000 30.170 4.280 ;
        RECT 31.010 4.000 33.480 4.280 ;
      LAYER met3 ;
        RECT 4.400 43.160 30.165 44.025 ;
        RECT 4.000 40.480 30.165 43.160 ;
        RECT 4.000 39.080 29.765 40.480 ;
        RECT 4.000 29.600 30.165 39.080 ;
        RECT 4.400 28.200 30.165 29.600 ;
        RECT 4.000 25.520 30.165 28.200 ;
        RECT 4.000 24.120 29.765 25.520 ;
        RECT 4.000 14.640 30.165 24.120 ;
        RECT 4.400 13.240 30.165 14.640 ;
        RECT 4.000 10.560 30.165 13.240 ;
        RECT 4.000 9.710 29.765 10.560 ;
      LAYER met4 ;
        RECT 8.575 10.640 25.590 43.760 ;
      LAYER met5 ;
        RECT 5.520 24.085 28.520 39.045 ;
  END
END dvsd_pe
END LIBRARY

