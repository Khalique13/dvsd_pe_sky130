magic
tech sky130A
magscale 1 2
timestamp 1634271523
<< viali >>
rect 2145 7497 2179 7531
rect 1409 7429 1443 7463
rect 1593 7429 1627 7463
rect 2881 7361 2915 7395
rect 3157 7361 3191 7395
rect 4537 7361 4571 7395
rect 4813 7361 4847 7395
rect 5273 7361 5307 7395
rect 7021 7361 7055 7395
rect 7665 7361 7699 7395
rect 3801 7157 3835 7191
rect 5457 7157 5491 7191
rect 6837 7157 6871 7191
rect 7481 7157 7515 7191
rect 3893 6953 3927 6987
rect 2697 6817 2731 6851
rect 4353 6817 4387 6851
rect 1409 6749 1443 6783
rect 2881 6749 2915 6783
rect 3893 6749 3927 6783
rect 4077 6749 4111 6783
rect 4169 6749 4203 6783
rect 4445 6749 4479 6783
rect 4997 6749 5031 6783
rect 5089 6749 5123 6783
rect 7941 6681 7975 6715
rect 1593 6613 1627 6647
rect 8033 6613 8067 6647
rect 3065 6409 3099 6443
rect 4077 6409 4111 6443
rect 4445 6341 4479 6375
rect 2973 6273 3007 6307
rect 3249 6273 3283 6307
rect 4261 6273 4295 6307
rect 4353 6273 4387 6307
rect 4629 6273 4663 6307
rect 4721 6273 4755 6307
rect 3249 6137 3283 6171
rect 3065 5865 3099 5899
rect 4445 5729 4479 5763
rect 5549 5729 5583 5763
rect 2973 5661 3007 5695
rect 4353 5661 4387 5695
rect 4721 5661 4755 5695
rect 4813 5661 4847 5695
rect 5457 5661 5491 5695
rect 5641 5661 5675 5695
rect 4997 5593 5031 5627
rect 4537 5525 4571 5559
rect 2605 5321 2639 5355
rect 3801 5321 3835 5355
rect 4537 5321 4571 5355
rect 6469 5321 6503 5355
rect 2237 5253 2271 5287
rect 2421 5185 2455 5219
rect 2513 5185 2547 5219
rect 3433 5185 3467 5219
rect 3617 5185 3651 5219
rect 4629 5185 4663 5219
rect 5273 5185 5307 5219
rect 5457 5185 5491 5219
rect 5549 5185 5583 5219
rect 6561 5185 6595 5219
rect 2789 5117 2823 5151
rect 5365 4981 5399 5015
rect 5733 4981 5767 5015
rect 4353 4777 4387 4811
rect 5273 4777 5307 4811
rect 4261 4573 4295 4607
rect 5457 4573 5491 4607
rect 4813 4097 4847 4131
rect 5089 4097 5123 4131
rect 7021 4097 7055 4131
rect 5825 3893 5859 3927
rect 7113 3893 7147 3927
rect 1593 3689 1627 3723
rect 1409 3485 1443 3519
rect 7941 3485 7975 3519
rect 8033 3349 8067 3383
rect 7941 3145 7975 3179
rect 8125 3009 8159 3043
rect 1593 2601 1627 2635
rect 2697 2601 2731 2635
rect 5089 2601 5123 2635
rect 1409 2397 1443 2431
rect 2513 2397 2547 2431
rect 4905 2397 4939 2431
rect 7481 2397 7515 2431
rect 7297 2329 7331 2363
<< metal1 >>
rect 1104 7642 8832 7664
rect 1104 7590 3547 7642
rect 3599 7590 3611 7642
rect 3663 7590 3675 7642
rect 3727 7590 3739 7642
rect 3791 7590 3803 7642
rect 3855 7590 6144 7642
rect 6196 7590 6208 7642
rect 6260 7590 6272 7642
rect 6324 7590 6336 7642
rect 6388 7590 6400 7642
rect 6452 7590 8832 7642
rect 1104 7568 8832 7590
rect 2133 7531 2191 7537
rect 2133 7497 2145 7531
rect 2179 7497 2191 7531
rect 2133 7491 2191 7497
rect 198 7420 204 7472
rect 256 7460 262 7472
rect 1397 7463 1455 7469
rect 1397 7460 1409 7463
rect 256 7432 1409 7460
rect 256 7420 262 7432
rect 1397 7429 1409 7432
rect 1443 7429 1455 7463
rect 1397 7423 1455 7429
rect 1581 7463 1639 7469
rect 1581 7429 1593 7463
rect 1627 7460 1639 7463
rect 2148 7460 2176 7491
rect 4154 7460 4160 7472
rect 1627 7432 2176 7460
rect 3160 7432 4160 7460
rect 1627 7429 1639 7432
rect 1581 7423 1639 7429
rect 2866 7392 2872 7404
rect 2827 7364 2872 7392
rect 2866 7352 2872 7364
rect 2924 7352 2930 7404
rect 3160 7401 3188 7432
rect 4154 7420 4160 7432
rect 4212 7460 4218 7472
rect 9766 7460 9772 7472
rect 4212 7432 4844 7460
rect 4212 7420 4218 7432
rect 3145 7395 3203 7401
rect 3145 7361 3157 7395
rect 3191 7361 3203 7395
rect 4522 7392 4528 7404
rect 4483 7364 4528 7392
rect 3145 7355 3203 7361
rect 4522 7352 4528 7364
rect 4580 7352 4586 7404
rect 4816 7401 4844 7432
rect 7024 7432 9772 7460
rect 4801 7395 4859 7401
rect 4801 7361 4813 7395
rect 4847 7361 4859 7395
rect 4801 7355 4859 7361
rect 4982 7352 4988 7404
rect 5040 7392 5046 7404
rect 7024 7401 7052 7432
rect 9766 7420 9772 7432
rect 9824 7420 9830 7472
rect 5261 7395 5319 7401
rect 5261 7392 5273 7395
rect 5040 7364 5273 7392
rect 5040 7352 5046 7364
rect 5261 7361 5273 7364
rect 5307 7361 5319 7395
rect 5261 7355 5319 7361
rect 7009 7395 7067 7401
rect 7009 7361 7021 7395
rect 7055 7361 7067 7395
rect 7009 7355 7067 7361
rect 7374 7352 7380 7404
rect 7432 7392 7438 7404
rect 7653 7395 7711 7401
rect 7653 7392 7665 7395
rect 7432 7364 7665 7392
rect 7432 7352 7438 7364
rect 7653 7361 7665 7364
rect 7699 7361 7711 7395
rect 7653 7355 7711 7361
rect 3786 7188 3792 7200
rect 3747 7160 3792 7188
rect 3786 7148 3792 7160
rect 3844 7148 3850 7200
rect 5442 7188 5448 7200
rect 5403 7160 5448 7188
rect 5442 7148 5448 7160
rect 5500 7148 5506 7200
rect 6822 7188 6828 7200
rect 6783 7160 6828 7188
rect 6822 7148 6828 7160
rect 6880 7148 6886 7200
rect 6914 7148 6920 7200
rect 6972 7188 6978 7200
rect 7469 7191 7527 7197
rect 7469 7188 7481 7191
rect 6972 7160 7481 7188
rect 6972 7148 6978 7160
rect 7469 7157 7481 7160
rect 7515 7157 7527 7191
rect 7469 7151 7527 7157
rect 1104 7098 8832 7120
rect 1104 7046 2248 7098
rect 2300 7046 2312 7098
rect 2364 7046 2376 7098
rect 2428 7046 2440 7098
rect 2492 7046 2504 7098
rect 2556 7046 4846 7098
rect 4898 7046 4910 7098
rect 4962 7046 4974 7098
rect 5026 7046 5038 7098
rect 5090 7046 5102 7098
rect 5154 7046 7443 7098
rect 7495 7046 7507 7098
rect 7559 7046 7571 7098
rect 7623 7046 7635 7098
rect 7687 7046 7699 7098
rect 7751 7046 8832 7098
rect 1104 7024 8832 7046
rect 2866 6944 2872 6996
rect 2924 6984 2930 6996
rect 3881 6987 3939 6993
rect 3881 6984 3893 6987
rect 2924 6956 3893 6984
rect 2924 6944 2930 6956
rect 3881 6953 3893 6956
rect 3927 6953 3939 6987
rect 3881 6947 3939 6953
rect 2590 6808 2596 6860
rect 2648 6848 2654 6860
rect 2685 6851 2743 6857
rect 2685 6848 2697 6851
rect 2648 6820 2697 6848
rect 2648 6808 2654 6820
rect 2685 6817 2697 6820
rect 2731 6817 2743 6851
rect 4246 6848 4252 6860
rect 2685 6811 2743 6817
rect 3896 6820 4252 6848
rect 1394 6780 1400 6792
rect 1355 6752 1400 6780
rect 1394 6740 1400 6752
rect 1452 6740 1458 6792
rect 2869 6783 2927 6789
rect 2869 6749 2881 6783
rect 2915 6780 2927 6783
rect 3786 6780 3792 6792
rect 2915 6752 3792 6780
rect 2915 6749 2927 6752
rect 2869 6743 2927 6749
rect 3786 6740 3792 6752
rect 3844 6740 3850 6792
rect 3896 6789 3924 6820
rect 4246 6808 4252 6820
rect 4304 6808 4310 6860
rect 4341 6851 4399 6857
rect 4341 6817 4353 6851
rect 4387 6848 4399 6851
rect 5534 6848 5540 6860
rect 4387 6820 5540 6848
rect 4387 6817 4399 6820
rect 4341 6811 4399 6817
rect 5534 6808 5540 6820
rect 5592 6848 5598 6860
rect 6822 6848 6828 6860
rect 5592 6820 6828 6848
rect 5592 6808 5598 6820
rect 6822 6808 6828 6820
rect 6880 6808 6886 6860
rect 3881 6783 3939 6789
rect 3881 6749 3893 6783
rect 3927 6749 3939 6783
rect 3881 6743 3939 6749
rect 4065 6783 4123 6789
rect 4065 6749 4077 6783
rect 4111 6749 4123 6783
rect 4065 6743 4123 6749
rect 1578 6644 1584 6656
rect 1539 6616 1584 6644
rect 1578 6604 1584 6616
rect 1636 6604 1642 6656
rect 4080 6644 4108 6743
rect 4154 6740 4160 6792
rect 4212 6780 4218 6792
rect 4430 6780 4436 6792
rect 4212 6752 4257 6780
rect 4343 6752 4436 6780
rect 4212 6740 4218 6752
rect 4430 6740 4436 6752
rect 4488 6780 4494 6792
rect 4985 6783 5043 6789
rect 4985 6780 4997 6783
rect 4488 6752 4997 6780
rect 4488 6740 4494 6752
rect 4985 6749 4997 6752
rect 5031 6749 5043 6783
rect 4985 6743 5043 6749
rect 5077 6783 5135 6789
rect 5077 6749 5089 6783
rect 5123 6780 5135 6783
rect 5442 6780 5448 6792
rect 5123 6752 5448 6780
rect 5123 6749 5135 6752
rect 5077 6743 5135 6749
rect 4246 6672 4252 6724
rect 4304 6712 4310 6724
rect 4614 6712 4620 6724
rect 4304 6684 4620 6712
rect 4304 6672 4310 6684
rect 4614 6672 4620 6684
rect 4672 6672 4678 6724
rect 4706 6672 4712 6724
rect 4764 6712 4770 6724
rect 5092 6712 5120 6743
rect 5442 6740 5448 6752
rect 5500 6740 5506 6792
rect 7926 6712 7932 6724
rect 4764 6684 5120 6712
rect 7887 6684 7932 6712
rect 4764 6672 4770 6684
rect 7926 6672 7932 6684
rect 7984 6672 7990 6724
rect 5166 6644 5172 6656
rect 4080 6616 5172 6644
rect 5166 6604 5172 6616
rect 5224 6604 5230 6656
rect 8018 6644 8024 6656
rect 7979 6616 8024 6644
rect 8018 6604 8024 6616
rect 8076 6604 8082 6656
rect 1104 6554 8832 6576
rect 1104 6502 3547 6554
rect 3599 6502 3611 6554
rect 3663 6502 3675 6554
rect 3727 6502 3739 6554
rect 3791 6502 3803 6554
rect 3855 6502 6144 6554
rect 6196 6502 6208 6554
rect 6260 6502 6272 6554
rect 6324 6502 6336 6554
rect 6388 6502 6400 6554
rect 6452 6502 8832 6554
rect 1104 6480 8832 6502
rect 1578 6400 1584 6452
rect 1636 6440 1642 6452
rect 2590 6440 2596 6452
rect 1636 6412 2596 6440
rect 1636 6400 1642 6412
rect 2590 6400 2596 6412
rect 2648 6440 2654 6452
rect 3053 6443 3111 6449
rect 3053 6440 3065 6443
rect 2648 6412 3065 6440
rect 2648 6400 2654 6412
rect 3053 6409 3065 6412
rect 3099 6409 3111 6443
rect 3053 6403 3111 6409
rect 4065 6443 4123 6449
rect 4065 6409 4077 6443
rect 4111 6440 4123 6443
rect 4522 6440 4528 6452
rect 4111 6412 4528 6440
rect 4111 6409 4123 6412
rect 4065 6403 4123 6409
rect 4522 6400 4528 6412
rect 4580 6400 4586 6452
rect 4430 6372 4436 6384
rect 4391 6344 4436 6372
rect 4430 6332 4436 6344
rect 4488 6332 4494 6384
rect 5534 6372 5540 6384
rect 4632 6344 5540 6372
rect 2958 6304 2964 6316
rect 2919 6276 2964 6304
rect 2958 6264 2964 6276
rect 3016 6264 3022 6316
rect 3237 6307 3295 6313
rect 3237 6273 3249 6307
rect 3283 6273 3295 6307
rect 4246 6304 4252 6316
rect 4207 6276 4252 6304
rect 3237 6267 3295 6273
rect 3252 6236 3280 6267
rect 4246 6264 4252 6276
rect 4304 6264 4310 6316
rect 4341 6307 4399 6313
rect 4341 6273 4353 6307
rect 4387 6273 4399 6307
rect 4341 6267 4399 6273
rect 3878 6236 3884 6248
rect 3252 6208 3884 6236
rect 3878 6196 3884 6208
rect 3936 6236 3942 6248
rect 4356 6236 4384 6267
rect 4522 6264 4528 6316
rect 4580 6304 4586 6316
rect 4632 6313 4660 6344
rect 5534 6332 5540 6344
rect 5592 6332 5598 6384
rect 4617 6307 4675 6313
rect 4617 6304 4629 6307
rect 4580 6276 4629 6304
rect 4580 6264 4586 6276
rect 4617 6273 4629 6276
rect 4663 6273 4675 6307
rect 4617 6267 4675 6273
rect 4709 6307 4767 6313
rect 4709 6273 4721 6307
rect 4755 6304 4767 6307
rect 5258 6304 5264 6316
rect 4755 6276 5264 6304
rect 4755 6273 4767 6276
rect 4709 6267 4767 6273
rect 5258 6264 5264 6276
rect 5316 6264 5322 6316
rect 5626 6236 5632 6248
rect 3936 6208 4292 6236
rect 4356 6208 5632 6236
rect 3936 6196 3942 6208
rect 3237 6171 3295 6177
rect 3237 6137 3249 6171
rect 3283 6168 3295 6171
rect 4154 6168 4160 6180
rect 3283 6140 4160 6168
rect 3283 6137 3295 6140
rect 3237 6131 3295 6137
rect 4154 6128 4160 6140
rect 4212 6128 4218 6180
rect 4264 6168 4292 6208
rect 5626 6196 5632 6208
rect 5684 6196 5690 6248
rect 6914 6168 6920 6180
rect 4264 6140 6920 6168
rect 6914 6128 6920 6140
rect 6972 6128 6978 6180
rect 1104 6010 8832 6032
rect 1104 5958 2248 6010
rect 2300 5958 2312 6010
rect 2364 5958 2376 6010
rect 2428 5958 2440 6010
rect 2492 5958 2504 6010
rect 2556 5958 4846 6010
rect 4898 5958 4910 6010
rect 4962 5958 4974 6010
rect 5026 5958 5038 6010
rect 5090 5958 5102 6010
rect 5154 5958 7443 6010
rect 7495 5958 7507 6010
rect 7559 5958 7571 6010
rect 7623 5958 7635 6010
rect 7687 5958 7699 6010
rect 7751 5958 8832 6010
rect 1104 5936 8832 5958
rect 2958 5856 2964 5908
rect 3016 5896 3022 5908
rect 3053 5899 3111 5905
rect 3053 5896 3065 5899
rect 3016 5868 3065 5896
rect 3016 5856 3022 5868
rect 3053 5865 3065 5868
rect 3099 5865 3111 5899
rect 3053 5859 3111 5865
rect 4433 5763 4491 5769
rect 4433 5729 4445 5763
rect 4479 5760 4491 5763
rect 5537 5763 5595 5769
rect 5537 5760 5549 5763
rect 4479 5732 5549 5760
rect 4479 5729 4491 5732
rect 4433 5723 4491 5729
rect 5537 5729 5549 5732
rect 5583 5729 5595 5763
rect 5537 5723 5595 5729
rect 2958 5692 2964 5704
rect 2919 5664 2964 5692
rect 2958 5652 2964 5664
rect 3016 5652 3022 5704
rect 4338 5692 4344 5704
rect 4299 5664 4344 5692
rect 4338 5652 4344 5664
rect 4396 5652 4402 5704
rect 4706 5692 4712 5704
rect 4667 5664 4712 5692
rect 4706 5652 4712 5664
rect 4764 5652 4770 5704
rect 4801 5695 4859 5701
rect 4801 5661 4813 5695
rect 4847 5661 4859 5695
rect 5445 5695 5503 5701
rect 5445 5692 5457 5695
rect 4801 5655 4859 5661
rect 4908 5664 5457 5692
rect 4430 5584 4436 5636
rect 4488 5624 4494 5636
rect 4816 5624 4844 5655
rect 4488 5596 4844 5624
rect 4488 5584 4494 5596
rect 4522 5556 4528 5568
rect 4483 5528 4528 5556
rect 4522 5516 4528 5528
rect 4580 5516 4586 5568
rect 4614 5516 4620 5568
rect 4672 5556 4678 5568
rect 4908 5556 4936 5664
rect 5445 5661 5457 5664
rect 5491 5661 5503 5695
rect 5626 5692 5632 5704
rect 5587 5664 5632 5692
rect 5445 5655 5503 5661
rect 5626 5652 5632 5664
rect 5684 5652 5690 5704
rect 4985 5627 5043 5633
rect 4985 5593 4997 5627
rect 5031 5624 5043 5627
rect 7006 5624 7012 5636
rect 5031 5596 7012 5624
rect 5031 5593 5043 5596
rect 4985 5587 5043 5593
rect 7006 5584 7012 5596
rect 7064 5624 7070 5636
rect 7926 5624 7932 5636
rect 7064 5596 7932 5624
rect 7064 5584 7070 5596
rect 7926 5584 7932 5596
rect 7984 5584 7990 5636
rect 4672 5528 4936 5556
rect 4672 5516 4678 5528
rect 1104 5466 8832 5488
rect 1104 5414 3547 5466
rect 3599 5414 3611 5466
rect 3663 5414 3675 5466
rect 3727 5414 3739 5466
rect 3791 5414 3803 5466
rect 3855 5414 6144 5466
rect 6196 5414 6208 5466
rect 6260 5414 6272 5466
rect 6324 5414 6336 5466
rect 6388 5414 6400 5466
rect 6452 5414 8832 5466
rect 1104 5392 8832 5414
rect 2590 5352 2596 5364
rect 2551 5324 2596 5352
rect 2590 5312 2596 5324
rect 2648 5312 2654 5364
rect 3789 5355 3847 5361
rect 3789 5321 3801 5355
rect 3835 5352 3847 5355
rect 4246 5352 4252 5364
rect 3835 5324 4252 5352
rect 3835 5321 3847 5324
rect 3789 5315 3847 5321
rect 4246 5312 4252 5324
rect 4304 5312 4310 5364
rect 4525 5355 4583 5361
rect 4525 5321 4537 5355
rect 4571 5352 4583 5355
rect 4614 5352 4620 5364
rect 4571 5324 4620 5352
rect 4571 5321 4583 5324
rect 4525 5315 4583 5321
rect 4614 5312 4620 5324
rect 4672 5312 4678 5364
rect 5626 5312 5632 5364
rect 5684 5352 5690 5364
rect 6457 5355 6515 5361
rect 6457 5352 6469 5355
rect 5684 5324 6469 5352
rect 5684 5312 5690 5324
rect 6457 5321 6469 5324
rect 6503 5321 6515 5355
rect 6457 5315 6515 5321
rect 2225 5287 2283 5293
rect 2225 5253 2237 5287
rect 2271 5284 2283 5287
rect 4338 5284 4344 5296
rect 2271 5256 4344 5284
rect 2271 5253 2283 5256
rect 2225 5247 2283 5253
rect 4338 5244 4344 5256
rect 4396 5244 4402 5296
rect 4706 5244 4712 5296
rect 4764 5284 4770 5296
rect 4764 5256 5580 5284
rect 4764 5244 4770 5256
rect 1578 5176 1584 5228
rect 1636 5216 1642 5228
rect 2409 5219 2467 5225
rect 2409 5216 2421 5219
rect 1636 5188 2421 5216
rect 1636 5176 1642 5188
rect 2409 5185 2421 5188
rect 2455 5185 2467 5219
rect 2409 5179 2467 5185
rect 2501 5219 2559 5225
rect 2501 5185 2513 5219
rect 2547 5216 2559 5219
rect 2958 5216 2964 5228
rect 2547 5188 2964 5216
rect 2547 5185 2559 5188
rect 2501 5179 2559 5185
rect 2130 5108 2136 5160
rect 2188 5148 2194 5160
rect 2516 5148 2544 5179
rect 2958 5176 2964 5188
rect 3016 5216 3022 5228
rect 3421 5219 3479 5225
rect 3421 5216 3433 5219
rect 3016 5188 3433 5216
rect 3016 5176 3022 5188
rect 3421 5185 3433 5188
rect 3467 5185 3479 5219
rect 3421 5179 3479 5185
rect 3605 5219 3663 5225
rect 3605 5185 3617 5219
rect 3651 5216 3663 5219
rect 3878 5216 3884 5228
rect 3651 5188 3884 5216
rect 3651 5185 3663 5188
rect 3605 5179 3663 5185
rect 2188 5120 2544 5148
rect 2777 5151 2835 5157
rect 2188 5108 2194 5120
rect 2777 5117 2789 5151
rect 2823 5148 2835 5151
rect 3620 5148 3648 5179
rect 3878 5176 3884 5188
rect 3936 5176 3942 5228
rect 4617 5219 4675 5225
rect 4617 5185 4629 5219
rect 4663 5216 4675 5219
rect 5258 5216 5264 5228
rect 4663 5188 5264 5216
rect 4663 5185 4675 5188
rect 4617 5179 4675 5185
rect 5258 5176 5264 5188
rect 5316 5176 5322 5228
rect 5442 5216 5448 5228
rect 5403 5188 5448 5216
rect 5442 5176 5448 5188
rect 5500 5176 5506 5228
rect 5552 5225 5580 5256
rect 5537 5219 5595 5225
rect 5537 5185 5549 5219
rect 5583 5185 5595 5219
rect 6546 5216 6552 5228
rect 6507 5188 6552 5216
rect 5537 5179 5595 5185
rect 6546 5176 6552 5188
rect 6604 5176 6610 5228
rect 2823 5120 3648 5148
rect 2823 5117 2835 5120
rect 2777 5111 2835 5117
rect 6546 5080 6552 5092
rect 5368 5052 6552 5080
rect 5368 5021 5396 5052
rect 6546 5040 6552 5052
rect 6604 5040 6610 5092
rect 5353 5015 5411 5021
rect 5353 4981 5365 5015
rect 5399 4981 5411 5015
rect 5353 4975 5411 4981
rect 5442 4972 5448 5024
rect 5500 5012 5506 5024
rect 5721 5015 5779 5021
rect 5721 5012 5733 5015
rect 5500 4984 5733 5012
rect 5500 4972 5506 4984
rect 5721 4981 5733 4984
rect 5767 4981 5779 5015
rect 5721 4975 5779 4981
rect 1104 4922 8832 4944
rect 1104 4870 2248 4922
rect 2300 4870 2312 4922
rect 2364 4870 2376 4922
rect 2428 4870 2440 4922
rect 2492 4870 2504 4922
rect 2556 4870 4846 4922
rect 4898 4870 4910 4922
rect 4962 4870 4974 4922
rect 5026 4870 5038 4922
rect 5090 4870 5102 4922
rect 5154 4870 7443 4922
rect 7495 4870 7507 4922
rect 7559 4870 7571 4922
rect 7623 4870 7635 4922
rect 7687 4870 7699 4922
rect 7751 4870 8832 4922
rect 1104 4848 8832 4870
rect 4341 4811 4399 4817
rect 4341 4777 4353 4811
rect 4387 4808 4399 4811
rect 4430 4808 4436 4820
rect 4387 4780 4436 4808
rect 4387 4777 4399 4780
rect 4341 4771 4399 4777
rect 4430 4768 4436 4780
rect 4488 4768 4494 4820
rect 5166 4768 5172 4820
rect 5224 4808 5230 4820
rect 5261 4811 5319 4817
rect 5261 4808 5273 4811
rect 5224 4780 5273 4808
rect 5224 4768 5230 4780
rect 5261 4777 5273 4780
rect 5307 4777 5319 4811
rect 5261 4771 5319 4777
rect 4246 4604 4252 4616
rect 4207 4576 4252 4604
rect 4246 4564 4252 4576
rect 4304 4564 4310 4616
rect 5442 4604 5448 4616
rect 5403 4576 5448 4604
rect 5442 4564 5448 4576
rect 5500 4564 5506 4616
rect 1104 4378 8832 4400
rect 1104 4326 3547 4378
rect 3599 4326 3611 4378
rect 3663 4326 3675 4378
rect 3727 4326 3739 4378
rect 3791 4326 3803 4378
rect 3855 4326 6144 4378
rect 6196 4326 6208 4378
rect 6260 4326 6272 4378
rect 6324 4326 6336 4378
rect 6388 4326 6400 4378
rect 6452 4326 8832 4378
rect 1104 4304 8832 4326
rect 4246 4088 4252 4140
rect 4304 4128 4310 4140
rect 4801 4131 4859 4137
rect 4801 4128 4813 4131
rect 4304 4100 4813 4128
rect 4304 4088 4310 4100
rect 4801 4097 4813 4100
rect 4847 4097 4859 4131
rect 4801 4091 4859 4097
rect 5077 4131 5135 4137
rect 5077 4097 5089 4131
rect 5123 4128 5135 4131
rect 5166 4128 5172 4140
rect 5123 4100 5172 4128
rect 5123 4097 5135 4100
rect 5077 4091 5135 4097
rect 5166 4088 5172 4100
rect 5224 4088 5230 4140
rect 7006 4128 7012 4140
rect 6967 4100 7012 4128
rect 7006 4088 7012 4100
rect 7064 4088 7070 4140
rect 5810 3924 5816 3936
rect 5771 3896 5816 3924
rect 5810 3884 5816 3896
rect 5868 3884 5874 3936
rect 7098 3924 7104 3936
rect 7059 3896 7104 3924
rect 7098 3884 7104 3896
rect 7156 3884 7162 3936
rect 1104 3834 8832 3856
rect 1104 3782 2248 3834
rect 2300 3782 2312 3834
rect 2364 3782 2376 3834
rect 2428 3782 2440 3834
rect 2492 3782 2504 3834
rect 2556 3782 4846 3834
rect 4898 3782 4910 3834
rect 4962 3782 4974 3834
rect 5026 3782 5038 3834
rect 5090 3782 5102 3834
rect 5154 3782 7443 3834
rect 7495 3782 7507 3834
rect 7559 3782 7571 3834
rect 7623 3782 7635 3834
rect 7687 3782 7699 3834
rect 7751 3782 8832 3834
rect 1104 3760 8832 3782
rect 1578 3720 1584 3732
rect 1539 3692 1584 3720
rect 1578 3680 1584 3692
rect 1636 3680 1642 3732
rect 1394 3516 1400 3528
rect 1355 3488 1400 3516
rect 1394 3476 1400 3488
rect 1452 3476 1458 3528
rect 5810 3476 5816 3528
rect 5868 3516 5874 3528
rect 7929 3519 7987 3525
rect 7929 3516 7941 3519
rect 5868 3488 7941 3516
rect 5868 3476 5874 3488
rect 7929 3485 7941 3488
rect 7975 3485 7987 3519
rect 7929 3479 7987 3485
rect 8018 3380 8024 3392
rect 7979 3352 8024 3380
rect 8018 3340 8024 3352
rect 8076 3340 8082 3392
rect 1104 3290 8832 3312
rect 1104 3238 3547 3290
rect 3599 3238 3611 3290
rect 3663 3238 3675 3290
rect 3727 3238 3739 3290
rect 3791 3238 3803 3290
rect 3855 3238 6144 3290
rect 6196 3238 6208 3290
rect 6260 3238 6272 3290
rect 6324 3238 6336 3290
rect 6388 3238 6400 3290
rect 6452 3238 8832 3290
rect 1104 3216 8832 3238
rect 6546 3136 6552 3188
rect 6604 3176 6610 3188
rect 7929 3179 7987 3185
rect 7929 3176 7941 3179
rect 6604 3148 7941 3176
rect 6604 3136 6610 3148
rect 7929 3145 7941 3148
rect 7975 3145 7987 3179
rect 7929 3139 7987 3145
rect 8113 3043 8171 3049
rect 8113 3009 8125 3043
rect 8159 3040 8171 3043
rect 9582 3040 9588 3052
rect 8159 3012 9588 3040
rect 8159 3009 8171 3012
rect 8113 3003 8171 3009
rect 9582 3000 9588 3012
rect 9640 3000 9646 3052
rect 1104 2746 8832 2768
rect 1104 2694 2248 2746
rect 2300 2694 2312 2746
rect 2364 2694 2376 2746
rect 2428 2694 2440 2746
rect 2492 2694 2504 2746
rect 2556 2694 4846 2746
rect 4898 2694 4910 2746
rect 4962 2694 4974 2746
rect 5026 2694 5038 2746
rect 5090 2694 5102 2746
rect 5154 2694 7443 2746
rect 7495 2694 7507 2746
rect 7559 2694 7571 2746
rect 7623 2694 7635 2746
rect 7687 2694 7699 2746
rect 7751 2694 8832 2746
rect 1104 2672 8832 2694
rect 1581 2635 1639 2641
rect 1581 2601 1593 2635
rect 1627 2632 1639 2635
rect 2130 2632 2136 2644
rect 1627 2604 2136 2632
rect 1627 2601 1639 2604
rect 1581 2595 1639 2601
rect 2130 2592 2136 2604
rect 2188 2592 2194 2644
rect 2685 2635 2743 2641
rect 2685 2601 2697 2635
rect 2731 2632 2743 2635
rect 4246 2632 4252 2644
rect 2731 2604 4252 2632
rect 2731 2601 2743 2604
rect 2685 2595 2743 2601
rect 4246 2592 4252 2604
rect 4304 2592 4310 2644
rect 5077 2635 5135 2641
rect 5077 2601 5089 2635
rect 5123 2632 5135 2635
rect 5258 2632 5264 2644
rect 5123 2604 5264 2632
rect 5123 2601 5135 2604
rect 5077 2595 5135 2601
rect 5258 2592 5264 2604
rect 5316 2592 5322 2644
rect 14 2388 20 2440
rect 72 2428 78 2440
rect 1397 2431 1455 2437
rect 1397 2428 1409 2431
rect 72 2400 1409 2428
rect 72 2388 78 2400
rect 1397 2397 1409 2400
rect 1443 2397 1455 2431
rect 1397 2391 1455 2397
rect 2406 2388 2412 2440
rect 2464 2428 2470 2440
rect 2501 2431 2559 2437
rect 2501 2428 2513 2431
rect 2464 2400 2513 2428
rect 2464 2388 2470 2400
rect 2501 2397 2513 2400
rect 2547 2397 2559 2431
rect 2501 2391 2559 2397
rect 4798 2388 4804 2440
rect 4856 2428 4862 2440
rect 4893 2431 4951 2437
rect 4893 2428 4905 2431
rect 4856 2400 4905 2428
rect 4856 2388 4862 2400
rect 4893 2397 4905 2400
rect 4939 2397 4951 2431
rect 4893 2391 4951 2397
rect 7098 2388 7104 2440
rect 7156 2428 7162 2440
rect 7469 2431 7527 2437
rect 7469 2428 7481 2431
rect 7156 2400 7481 2428
rect 7156 2388 7162 2400
rect 7469 2397 7481 2400
rect 7515 2397 7527 2431
rect 7469 2391 7527 2397
rect 7190 2320 7196 2372
rect 7248 2360 7254 2372
rect 7285 2363 7343 2369
rect 7285 2360 7297 2363
rect 7248 2332 7297 2360
rect 7248 2320 7254 2332
rect 7285 2329 7297 2332
rect 7331 2329 7343 2363
rect 7285 2323 7343 2329
rect 1104 2202 8832 2224
rect 1104 2150 3547 2202
rect 3599 2150 3611 2202
rect 3663 2150 3675 2202
rect 3727 2150 3739 2202
rect 3791 2150 3803 2202
rect 3855 2150 6144 2202
rect 6196 2150 6208 2202
rect 6260 2150 6272 2202
rect 6324 2150 6336 2202
rect 6388 2150 6400 2202
rect 6452 2150 8832 2202
rect 1104 2128 8832 2150
<< via1 >>
rect 3547 7590 3599 7642
rect 3611 7590 3663 7642
rect 3675 7590 3727 7642
rect 3739 7590 3791 7642
rect 3803 7590 3855 7642
rect 6144 7590 6196 7642
rect 6208 7590 6260 7642
rect 6272 7590 6324 7642
rect 6336 7590 6388 7642
rect 6400 7590 6452 7642
rect 204 7420 256 7472
rect 2872 7395 2924 7404
rect 2872 7361 2881 7395
rect 2881 7361 2915 7395
rect 2915 7361 2924 7395
rect 2872 7352 2924 7361
rect 4160 7420 4212 7472
rect 4528 7395 4580 7404
rect 4528 7361 4537 7395
rect 4537 7361 4571 7395
rect 4571 7361 4580 7395
rect 4528 7352 4580 7361
rect 4988 7352 5040 7404
rect 9772 7420 9824 7472
rect 7380 7352 7432 7404
rect 3792 7191 3844 7200
rect 3792 7157 3801 7191
rect 3801 7157 3835 7191
rect 3835 7157 3844 7191
rect 3792 7148 3844 7157
rect 5448 7191 5500 7200
rect 5448 7157 5457 7191
rect 5457 7157 5491 7191
rect 5491 7157 5500 7191
rect 5448 7148 5500 7157
rect 6828 7191 6880 7200
rect 6828 7157 6837 7191
rect 6837 7157 6871 7191
rect 6871 7157 6880 7191
rect 6828 7148 6880 7157
rect 6920 7148 6972 7200
rect 2248 7046 2300 7098
rect 2312 7046 2364 7098
rect 2376 7046 2428 7098
rect 2440 7046 2492 7098
rect 2504 7046 2556 7098
rect 4846 7046 4898 7098
rect 4910 7046 4962 7098
rect 4974 7046 5026 7098
rect 5038 7046 5090 7098
rect 5102 7046 5154 7098
rect 7443 7046 7495 7098
rect 7507 7046 7559 7098
rect 7571 7046 7623 7098
rect 7635 7046 7687 7098
rect 7699 7046 7751 7098
rect 2872 6944 2924 6996
rect 2596 6808 2648 6860
rect 1400 6783 1452 6792
rect 1400 6749 1409 6783
rect 1409 6749 1443 6783
rect 1443 6749 1452 6783
rect 1400 6740 1452 6749
rect 3792 6740 3844 6792
rect 4252 6808 4304 6860
rect 5540 6808 5592 6860
rect 6828 6808 6880 6860
rect 1584 6647 1636 6656
rect 1584 6613 1593 6647
rect 1593 6613 1627 6647
rect 1627 6613 1636 6647
rect 1584 6604 1636 6613
rect 4160 6783 4212 6792
rect 4160 6749 4169 6783
rect 4169 6749 4203 6783
rect 4203 6749 4212 6783
rect 4436 6783 4488 6792
rect 4160 6740 4212 6749
rect 4436 6749 4445 6783
rect 4445 6749 4479 6783
rect 4479 6749 4488 6783
rect 4436 6740 4488 6749
rect 4252 6672 4304 6724
rect 4620 6672 4672 6724
rect 4712 6672 4764 6724
rect 5448 6740 5500 6792
rect 7932 6715 7984 6724
rect 7932 6681 7941 6715
rect 7941 6681 7975 6715
rect 7975 6681 7984 6715
rect 7932 6672 7984 6681
rect 5172 6604 5224 6656
rect 8024 6647 8076 6656
rect 8024 6613 8033 6647
rect 8033 6613 8067 6647
rect 8067 6613 8076 6647
rect 8024 6604 8076 6613
rect 3547 6502 3599 6554
rect 3611 6502 3663 6554
rect 3675 6502 3727 6554
rect 3739 6502 3791 6554
rect 3803 6502 3855 6554
rect 6144 6502 6196 6554
rect 6208 6502 6260 6554
rect 6272 6502 6324 6554
rect 6336 6502 6388 6554
rect 6400 6502 6452 6554
rect 1584 6400 1636 6452
rect 2596 6400 2648 6452
rect 4528 6400 4580 6452
rect 4436 6375 4488 6384
rect 4436 6341 4445 6375
rect 4445 6341 4479 6375
rect 4479 6341 4488 6375
rect 4436 6332 4488 6341
rect 2964 6307 3016 6316
rect 2964 6273 2973 6307
rect 2973 6273 3007 6307
rect 3007 6273 3016 6307
rect 2964 6264 3016 6273
rect 4252 6307 4304 6316
rect 4252 6273 4261 6307
rect 4261 6273 4295 6307
rect 4295 6273 4304 6307
rect 4252 6264 4304 6273
rect 3884 6196 3936 6248
rect 4528 6264 4580 6316
rect 5540 6332 5592 6384
rect 5264 6264 5316 6316
rect 4160 6128 4212 6180
rect 5632 6196 5684 6248
rect 6920 6128 6972 6180
rect 2248 5958 2300 6010
rect 2312 5958 2364 6010
rect 2376 5958 2428 6010
rect 2440 5958 2492 6010
rect 2504 5958 2556 6010
rect 4846 5958 4898 6010
rect 4910 5958 4962 6010
rect 4974 5958 5026 6010
rect 5038 5958 5090 6010
rect 5102 5958 5154 6010
rect 7443 5958 7495 6010
rect 7507 5958 7559 6010
rect 7571 5958 7623 6010
rect 7635 5958 7687 6010
rect 7699 5958 7751 6010
rect 2964 5856 3016 5908
rect 2964 5695 3016 5704
rect 2964 5661 2973 5695
rect 2973 5661 3007 5695
rect 3007 5661 3016 5695
rect 2964 5652 3016 5661
rect 4344 5695 4396 5704
rect 4344 5661 4353 5695
rect 4353 5661 4387 5695
rect 4387 5661 4396 5695
rect 4344 5652 4396 5661
rect 4712 5695 4764 5704
rect 4712 5661 4721 5695
rect 4721 5661 4755 5695
rect 4755 5661 4764 5695
rect 4712 5652 4764 5661
rect 4436 5584 4488 5636
rect 4528 5559 4580 5568
rect 4528 5525 4537 5559
rect 4537 5525 4571 5559
rect 4571 5525 4580 5559
rect 4528 5516 4580 5525
rect 4620 5516 4672 5568
rect 5632 5695 5684 5704
rect 5632 5661 5641 5695
rect 5641 5661 5675 5695
rect 5675 5661 5684 5695
rect 5632 5652 5684 5661
rect 7012 5584 7064 5636
rect 7932 5584 7984 5636
rect 3547 5414 3599 5466
rect 3611 5414 3663 5466
rect 3675 5414 3727 5466
rect 3739 5414 3791 5466
rect 3803 5414 3855 5466
rect 6144 5414 6196 5466
rect 6208 5414 6260 5466
rect 6272 5414 6324 5466
rect 6336 5414 6388 5466
rect 6400 5414 6452 5466
rect 2596 5355 2648 5364
rect 2596 5321 2605 5355
rect 2605 5321 2639 5355
rect 2639 5321 2648 5355
rect 2596 5312 2648 5321
rect 4252 5312 4304 5364
rect 4620 5312 4672 5364
rect 5632 5312 5684 5364
rect 4344 5244 4396 5296
rect 4712 5244 4764 5296
rect 1584 5176 1636 5228
rect 2136 5108 2188 5160
rect 2964 5176 3016 5228
rect 3884 5176 3936 5228
rect 5264 5219 5316 5228
rect 5264 5185 5273 5219
rect 5273 5185 5307 5219
rect 5307 5185 5316 5219
rect 5264 5176 5316 5185
rect 5448 5219 5500 5228
rect 5448 5185 5457 5219
rect 5457 5185 5491 5219
rect 5491 5185 5500 5219
rect 5448 5176 5500 5185
rect 6552 5219 6604 5228
rect 6552 5185 6561 5219
rect 6561 5185 6595 5219
rect 6595 5185 6604 5219
rect 6552 5176 6604 5185
rect 6552 5040 6604 5092
rect 5448 4972 5500 5024
rect 2248 4870 2300 4922
rect 2312 4870 2364 4922
rect 2376 4870 2428 4922
rect 2440 4870 2492 4922
rect 2504 4870 2556 4922
rect 4846 4870 4898 4922
rect 4910 4870 4962 4922
rect 4974 4870 5026 4922
rect 5038 4870 5090 4922
rect 5102 4870 5154 4922
rect 7443 4870 7495 4922
rect 7507 4870 7559 4922
rect 7571 4870 7623 4922
rect 7635 4870 7687 4922
rect 7699 4870 7751 4922
rect 4436 4768 4488 4820
rect 5172 4768 5224 4820
rect 4252 4607 4304 4616
rect 4252 4573 4261 4607
rect 4261 4573 4295 4607
rect 4295 4573 4304 4607
rect 4252 4564 4304 4573
rect 5448 4607 5500 4616
rect 5448 4573 5457 4607
rect 5457 4573 5491 4607
rect 5491 4573 5500 4607
rect 5448 4564 5500 4573
rect 3547 4326 3599 4378
rect 3611 4326 3663 4378
rect 3675 4326 3727 4378
rect 3739 4326 3791 4378
rect 3803 4326 3855 4378
rect 6144 4326 6196 4378
rect 6208 4326 6260 4378
rect 6272 4326 6324 4378
rect 6336 4326 6388 4378
rect 6400 4326 6452 4378
rect 4252 4088 4304 4140
rect 5172 4088 5224 4140
rect 7012 4131 7064 4140
rect 7012 4097 7021 4131
rect 7021 4097 7055 4131
rect 7055 4097 7064 4131
rect 7012 4088 7064 4097
rect 5816 3927 5868 3936
rect 5816 3893 5825 3927
rect 5825 3893 5859 3927
rect 5859 3893 5868 3927
rect 5816 3884 5868 3893
rect 7104 3927 7156 3936
rect 7104 3893 7113 3927
rect 7113 3893 7147 3927
rect 7147 3893 7156 3927
rect 7104 3884 7156 3893
rect 2248 3782 2300 3834
rect 2312 3782 2364 3834
rect 2376 3782 2428 3834
rect 2440 3782 2492 3834
rect 2504 3782 2556 3834
rect 4846 3782 4898 3834
rect 4910 3782 4962 3834
rect 4974 3782 5026 3834
rect 5038 3782 5090 3834
rect 5102 3782 5154 3834
rect 7443 3782 7495 3834
rect 7507 3782 7559 3834
rect 7571 3782 7623 3834
rect 7635 3782 7687 3834
rect 7699 3782 7751 3834
rect 1584 3723 1636 3732
rect 1584 3689 1593 3723
rect 1593 3689 1627 3723
rect 1627 3689 1636 3723
rect 1584 3680 1636 3689
rect 1400 3519 1452 3528
rect 1400 3485 1409 3519
rect 1409 3485 1443 3519
rect 1443 3485 1452 3519
rect 1400 3476 1452 3485
rect 5816 3476 5868 3528
rect 8024 3383 8076 3392
rect 8024 3349 8033 3383
rect 8033 3349 8067 3383
rect 8067 3349 8076 3383
rect 8024 3340 8076 3349
rect 3547 3238 3599 3290
rect 3611 3238 3663 3290
rect 3675 3238 3727 3290
rect 3739 3238 3791 3290
rect 3803 3238 3855 3290
rect 6144 3238 6196 3290
rect 6208 3238 6260 3290
rect 6272 3238 6324 3290
rect 6336 3238 6388 3290
rect 6400 3238 6452 3290
rect 6552 3136 6604 3188
rect 9588 3000 9640 3052
rect 2248 2694 2300 2746
rect 2312 2694 2364 2746
rect 2376 2694 2428 2746
rect 2440 2694 2492 2746
rect 2504 2694 2556 2746
rect 4846 2694 4898 2746
rect 4910 2694 4962 2746
rect 4974 2694 5026 2746
rect 5038 2694 5090 2746
rect 5102 2694 5154 2746
rect 7443 2694 7495 2746
rect 7507 2694 7559 2746
rect 7571 2694 7623 2746
rect 7635 2694 7687 2746
rect 7699 2694 7751 2746
rect 2136 2592 2188 2644
rect 4252 2592 4304 2644
rect 5264 2592 5316 2644
rect 20 2388 72 2440
rect 2412 2388 2464 2440
rect 4804 2388 4856 2440
rect 7104 2388 7156 2440
rect 7196 2320 7248 2372
rect 3547 2150 3599 2202
rect 3611 2150 3663 2202
rect 3675 2150 3727 2202
rect 3739 2150 3791 2202
rect 3803 2150 3855 2202
rect 6144 2150 6196 2202
rect 6208 2150 6260 2202
rect 6272 2150 6324 2202
rect 6336 2150 6388 2202
rect 6400 2150 6452 2202
<< metal2 >>
rect 202 9200 258 10000
rect 2594 9200 2650 10000
rect 4986 9200 5042 10000
rect 7378 9200 7434 10000
rect 9770 9200 9826 10000
rect 216 7478 244 9200
rect 204 7472 256 7478
rect 204 7414 256 7420
rect 2248 7100 2556 7120
rect 2248 7098 2254 7100
rect 2310 7098 2334 7100
rect 2390 7098 2414 7100
rect 2470 7098 2494 7100
rect 2550 7098 2556 7100
rect 2310 7046 2312 7098
rect 2492 7046 2494 7098
rect 2248 7044 2254 7046
rect 2310 7044 2334 7046
rect 2390 7044 2414 7046
rect 2470 7044 2494 7046
rect 2550 7044 2556 7046
rect 2248 7024 2556 7044
rect 1398 6896 1454 6905
rect 2608 6866 2636 9200
rect 3547 7644 3855 7664
rect 3547 7642 3553 7644
rect 3609 7642 3633 7644
rect 3689 7642 3713 7644
rect 3769 7642 3793 7644
rect 3849 7642 3855 7644
rect 3609 7590 3611 7642
rect 3791 7590 3793 7642
rect 3547 7588 3553 7590
rect 3609 7588 3633 7590
rect 3689 7588 3713 7590
rect 3769 7588 3793 7590
rect 3849 7588 3855 7590
rect 3547 7568 3855 7588
rect 4160 7472 4212 7478
rect 4160 7414 4212 7420
rect 2872 7404 2924 7410
rect 2872 7346 2924 7352
rect 2884 7002 2912 7346
rect 3792 7200 3844 7206
rect 3792 7142 3844 7148
rect 2872 6996 2924 7002
rect 2872 6938 2924 6944
rect 1398 6831 1454 6840
rect 2596 6860 2648 6866
rect 1412 6798 1440 6831
rect 2596 6802 2648 6808
rect 3804 6798 3832 7142
rect 4172 6882 4200 7414
rect 5000 7410 5028 9200
rect 6144 7644 6452 7664
rect 6144 7642 6150 7644
rect 6206 7642 6230 7644
rect 6286 7642 6310 7644
rect 6366 7642 6390 7644
rect 6446 7642 6452 7644
rect 6206 7590 6208 7642
rect 6388 7590 6390 7642
rect 6144 7588 6150 7590
rect 6206 7588 6230 7590
rect 6286 7588 6310 7590
rect 6366 7588 6390 7590
rect 6446 7588 6452 7590
rect 6144 7568 6452 7588
rect 7392 7410 7420 9200
rect 9784 7478 9812 9200
rect 9772 7472 9824 7478
rect 9772 7414 9824 7420
rect 4528 7404 4580 7410
rect 4528 7346 4580 7352
rect 4988 7404 5040 7410
rect 4988 7346 5040 7352
rect 7380 7404 7432 7410
rect 7380 7346 7432 7352
rect 4080 6854 4200 6882
rect 4252 6860 4304 6866
rect 1400 6792 1452 6798
rect 1400 6734 1452 6740
rect 3792 6792 3844 6798
rect 3792 6734 3844 6740
rect 1584 6656 1636 6662
rect 1584 6598 1636 6604
rect 1596 6458 1624 6598
rect 3547 6556 3855 6576
rect 3547 6554 3553 6556
rect 3609 6554 3633 6556
rect 3689 6554 3713 6556
rect 3769 6554 3793 6556
rect 3849 6554 3855 6556
rect 3609 6502 3611 6554
rect 3791 6502 3793 6554
rect 3547 6500 3553 6502
rect 3609 6500 3633 6502
rect 3689 6500 3713 6502
rect 3769 6500 3793 6502
rect 3849 6500 3855 6502
rect 3547 6480 3855 6500
rect 1584 6452 1636 6458
rect 1584 6394 1636 6400
rect 2596 6452 2648 6458
rect 2596 6394 2648 6400
rect 2248 6012 2556 6032
rect 2248 6010 2254 6012
rect 2310 6010 2334 6012
rect 2390 6010 2414 6012
rect 2470 6010 2494 6012
rect 2550 6010 2556 6012
rect 2310 5958 2312 6010
rect 2492 5958 2494 6010
rect 2248 5956 2254 5958
rect 2310 5956 2334 5958
rect 2390 5956 2414 5958
rect 2470 5956 2494 5958
rect 2550 5956 2556 5958
rect 2248 5936 2556 5956
rect 2608 5370 2636 6394
rect 2964 6316 3016 6322
rect 2964 6258 3016 6264
rect 2976 5914 3004 6258
rect 3884 6248 3936 6254
rect 3884 6190 3936 6196
rect 2964 5908 3016 5914
rect 2964 5850 3016 5856
rect 2964 5704 3016 5710
rect 2964 5646 3016 5652
rect 2596 5364 2648 5370
rect 2596 5306 2648 5312
rect 2976 5234 3004 5646
rect 3547 5468 3855 5488
rect 3547 5466 3553 5468
rect 3609 5466 3633 5468
rect 3689 5466 3713 5468
rect 3769 5466 3793 5468
rect 3849 5466 3855 5468
rect 3609 5414 3611 5466
rect 3791 5414 3793 5466
rect 3547 5412 3553 5414
rect 3609 5412 3633 5414
rect 3689 5412 3713 5414
rect 3769 5412 3793 5414
rect 3849 5412 3855 5414
rect 3547 5392 3855 5412
rect 3896 5234 3924 6190
rect 4080 6066 4108 6854
rect 4252 6802 4304 6808
rect 4160 6792 4212 6798
rect 4160 6734 4212 6740
rect 4172 6186 4200 6734
rect 4264 6730 4292 6802
rect 4436 6792 4488 6798
rect 4436 6734 4488 6740
rect 4252 6724 4304 6730
rect 4252 6666 4304 6672
rect 4448 6390 4476 6734
rect 4540 6458 4568 7346
rect 5448 7200 5500 7206
rect 5448 7142 5500 7148
rect 6828 7200 6880 7206
rect 6828 7142 6880 7148
rect 6920 7200 6972 7206
rect 6920 7142 6972 7148
rect 4846 7100 5154 7120
rect 4846 7098 4852 7100
rect 4908 7098 4932 7100
rect 4988 7098 5012 7100
rect 5068 7098 5092 7100
rect 5148 7098 5154 7100
rect 4908 7046 4910 7098
rect 5090 7046 5092 7098
rect 4846 7044 4852 7046
rect 4908 7044 4932 7046
rect 4988 7044 5012 7046
rect 5068 7044 5092 7046
rect 5148 7044 5154 7046
rect 4846 7024 5154 7044
rect 5460 6798 5488 7142
rect 6840 6866 6868 7142
rect 5540 6860 5592 6866
rect 5540 6802 5592 6808
rect 6828 6860 6880 6866
rect 6828 6802 6880 6808
rect 5448 6792 5500 6798
rect 5448 6734 5500 6740
rect 4620 6724 4672 6730
rect 4620 6666 4672 6672
rect 4712 6724 4764 6730
rect 4712 6666 4764 6672
rect 4528 6452 4580 6458
rect 4528 6394 4580 6400
rect 4436 6384 4488 6390
rect 4436 6326 4488 6332
rect 4252 6316 4304 6322
rect 4252 6258 4304 6264
rect 4528 6316 4580 6322
rect 4528 6258 4580 6264
rect 4160 6180 4212 6186
rect 4160 6122 4212 6128
rect 4080 6038 4200 6066
rect 1584 5228 1636 5234
rect 1584 5170 1636 5176
rect 2964 5228 3016 5234
rect 2964 5170 3016 5176
rect 3884 5228 3936 5234
rect 3884 5170 3936 5176
rect 1596 3738 1624 5170
rect 2136 5160 2188 5166
rect 2136 5102 2188 5108
rect 1584 3732 1636 3738
rect 1584 3674 1636 3680
rect 1400 3528 1452 3534
rect 1400 3470 1452 3476
rect 1412 3369 1440 3470
rect 1398 3360 1454 3369
rect 1398 3295 1454 3304
rect 2148 2650 2176 5102
rect 2248 4924 2556 4944
rect 2248 4922 2254 4924
rect 2310 4922 2334 4924
rect 2390 4922 2414 4924
rect 2470 4922 2494 4924
rect 2550 4922 2556 4924
rect 2310 4870 2312 4922
rect 2492 4870 2494 4922
rect 2248 4868 2254 4870
rect 2310 4868 2334 4870
rect 2390 4868 2414 4870
rect 2470 4868 2494 4870
rect 2550 4868 2556 4870
rect 2248 4848 2556 4868
rect 4172 4706 4200 6038
rect 4264 5370 4292 6258
rect 4344 5704 4396 5710
rect 4344 5646 4396 5652
rect 4252 5364 4304 5370
rect 4252 5306 4304 5312
rect 4356 5302 4384 5646
rect 4436 5636 4488 5642
rect 4436 5578 4488 5584
rect 4344 5296 4396 5302
rect 4344 5238 4396 5244
rect 4448 4826 4476 5578
rect 4540 5574 4568 6258
rect 4632 5574 4660 6666
rect 4724 5710 4752 6666
rect 5172 6656 5224 6662
rect 5172 6598 5224 6604
rect 4846 6012 5154 6032
rect 4846 6010 4852 6012
rect 4908 6010 4932 6012
rect 4988 6010 5012 6012
rect 5068 6010 5092 6012
rect 5148 6010 5154 6012
rect 4908 5958 4910 6010
rect 5090 5958 5092 6010
rect 4846 5956 4852 5958
rect 4908 5956 4932 5958
rect 4988 5956 5012 5958
rect 5068 5956 5092 5958
rect 5148 5956 5154 5958
rect 4846 5936 5154 5956
rect 4712 5704 4764 5710
rect 4712 5646 4764 5652
rect 4528 5568 4580 5574
rect 4528 5510 4580 5516
rect 4620 5568 4672 5574
rect 4620 5510 4672 5516
rect 4632 5370 4660 5510
rect 4620 5364 4672 5370
rect 4620 5306 4672 5312
rect 4724 5302 4752 5646
rect 4712 5296 4764 5302
rect 4712 5238 4764 5244
rect 4846 4924 5154 4944
rect 4846 4922 4852 4924
rect 4908 4922 4932 4924
rect 4988 4922 5012 4924
rect 5068 4922 5092 4924
rect 5148 4922 5154 4924
rect 4908 4870 4910 4922
rect 5090 4870 5092 4922
rect 4846 4868 4852 4870
rect 4908 4868 4932 4870
rect 4988 4868 5012 4870
rect 5068 4868 5092 4870
rect 5148 4868 5154 4870
rect 4846 4848 5154 4868
rect 5184 4826 5212 6598
rect 5552 6390 5580 6802
rect 6144 6556 6452 6576
rect 6144 6554 6150 6556
rect 6206 6554 6230 6556
rect 6286 6554 6310 6556
rect 6366 6554 6390 6556
rect 6446 6554 6452 6556
rect 6206 6502 6208 6554
rect 6388 6502 6390 6554
rect 6144 6500 6150 6502
rect 6206 6500 6230 6502
rect 6286 6500 6310 6502
rect 6366 6500 6390 6502
rect 6446 6500 6452 6502
rect 6144 6480 6452 6500
rect 5540 6384 5592 6390
rect 5540 6326 5592 6332
rect 5264 6316 5316 6322
rect 5264 6258 5316 6264
rect 5276 5234 5304 6258
rect 5552 5250 5580 6326
rect 5632 6248 5684 6254
rect 5632 6190 5684 6196
rect 5644 5710 5672 6190
rect 6932 6186 6960 7142
rect 7443 7100 7751 7120
rect 7443 7098 7449 7100
rect 7505 7098 7529 7100
rect 7585 7098 7609 7100
rect 7665 7098 7689 7100
rect 7745 7098 7751 7100
rect 7505 7046 7507 7098
rect 7687 7046 7689 7098
rect 7443 7044 7449 7046
rect 7505 7044 7529 7046
rect 7585 7044 7609 7046
rect 7665 7044 7689 7046
rect 7745 7044 7751 7046
rect 7443 7024 7751 7044
rect 7932 6724 7984 6730
rect 7932 6666 7984 6672
rect 6920 6180 6972 6186
rect 6920 6122 6972 6128
rect 7443 6012 7751 6032
rect 7443 6010 7449 6012
rect 7505 6010 7529 6012
rect 7585 6010 7609 6012
rect 7665 6010 7689 6012
rect 7745 6010 7751 6012
rect 7505 5958 7507 6010
rect 7687 5958 7689 6010
rect 7443 5956 7449 5958
rect 7505 5956 7529 5958
rect 7585 5956 7609 5958
rect 7665 5956 7689 5958
rect 7745 5956 7751 5958
rect 7443 5936 7751 5956
rect 5632 5704 5684 5710
rect 5632 5646 5684 5652
rect 5644 5370 5672 5646
rect 7944 5642 7972 6666
rect 8024 6656 8076 6662
rect 8022 6624 8024 6633
rect 8076 6624 8078 6633
rect 8022 6559 8078 6568
rect 7012 5636 7064 5642
rect 7012 5578 7064 5584
rect 7932 5636 7984 5642
rect 7932 5578 7984 5584
rect 6144 5468 6452 5488
rect 6144 5466 6150 5468
rect 6206 5466 6230 5468
rect 6286 5466 6310 5468
rect 6366 5466 6390 5468
rect 6446 5466 6452 5468
rect 6206 5414 6208 5466
rect 6388 5414 6390 5466
rect 6144 5412 6150 5414
rect 6206 5412 6230 5414
rect 6286 5412 6310 5414
rect 6366 5412 6390 5414
rect 6446 5412 6452 5414
rect 6144 5392 6452 5412
rect 5632 5364 5684 5370
rect 5632 5306 5684 5312
rect 5460 5234 5580 5250
rect 5264 5228 5316 5234
rect 5264 5170 5316 5176
rect 5448 5228 5580 5234
rect 5500 5222 5580 5228
rect 6552 5228 6604 5234
rect 5448 5170 5500 5176
rect 6552 5170 6604 5176
rect 4436 4820 4488 4826
rect 4436 4762 4488 4768
rect 5172 4820 5224 4826
rect 5172 4762 5224 4768
rect 4172 4678 4292 4706
rect 4264 4622 4292 4678
rect 4252 4616 4304 4622
rect 4252 4558 4304 4564
rect 3547 4380 3855 4400
rect 3547 4378 3553 4380
rect 3609 4378 3633 4380
rect 3689 4378 3713 4380
rect 3769 4378 3793 4380
rect 3849 4378 3855 4380
rect 3609 4326 3611 4378
rect 3791 4326 3793 4378
rect 3547 4324 3553 4326
rect 3609 4324 3633 4326
rect 3689 4324 3713 4326
rect 3769 4324 3793 4326
rect 3849 4324 3855 4326
rect 3547 4304 3855 4324
rect 4264 4146 4292 4558
rect 5184 4146 5212 4762
rect 4252 4140 4304 4146
rect 4252 4082 4304 4088
rect 5172 4140 5224 4146
rect 5172 4082 5224 4088
rect 2248 3836 2556 3856
rect 2248 3834 2254 3836
rect 2310 3834 2334 3836
rect 2390 3834 2414 3836
rect 2470 3834 2494 3836
rect 2550 3834 2556 3836
rect 2310 3782 2312 3834
rect 2492 3782 2494 3834
rect 2248 3780 2254 3782
rect 2310 3780 2334 3782
rect 2390 3780 2414 3782
rect 2470 3780 2494 3782
rect 2550 3780 2556 3782
rect 2248 3760 2556 3780
rect 3547 3292 3855 3312
rect 3547 3290 3553 3292
rect 3609 3290 3633 3292
rect 3689 3290 3713 3292
rect 3769 3290 3793 3292
rect 3849 3290 3855 3292
rect 3609 3238 3611 3290
rect 3791 3238 3793 3290
rect 3547 3236 3553 3238
rect 3609 3236 3633 3238
rect 3689 3236 3713 3238
rect 3769 3236 3793 3238
rect 3849 3236 3855 3238
rect 3547 3216 3855 3236
rect 2248 2748 2556 2768
rect 2248 2746 2254 2748
rect 2310 2746 2334 2748
rect 2390 2746 2414 2748
rect 2470 2746 2494 2748
rect 2550 2746 2556 2748
rect 2310 2694 2312 2746
rect 2492 2694 2494 2746
rect 2248 2692 2254 2694
rect 2310 2692 2334 2694
rect 2390 2692 2414 2694
rect 2470 2692 2494 2694
rect 2550 2692 2556 2694
rect 2248 2672 2556 2692
rect 4264 2650 4292 4082
rect 4846 3836 5154 3856
rect 4846 3834 4852 3836
rect 4908 3834 4932 3836
rect 4988 3834 5012 3836
rect 5068 3834 5092 3836
rect 5148 3834 5154 3836
rect 4908 3782 4910 3834
rect 5090 3782 5092 3834
rect 4846 3780 4852 3782
rect 4908 3780 4932 3782
rect 4988 3780 5012 3782
rect 5068 3780 5092 3782
rect 5148 3780 5154 3782
rect 4846 3760 5154 3780
rect 4846 2748 5154 2768
rect 4846 2746 4852 2748
rect 4908 2746 4932 2748
rect 4988 2746 5012 2748
rect 5068 2746 5092 2748
rect 5148 2746 5154 2748
rect 4908 2694 4910 2746
rect 5090 2694 5092 2746
rect 4846 2692 4852 2694
rect 4908 2692 4932 2694
rect 4988 2692 5012 2694
rect 5068 2692 5092 2694
rect 5148 2692 5154 2694
rect 4846 2672 5154 2692
rect 5276 2650 5304 5170
rect 6564 5098 6592 5170
rect 6552 5092 6604 5098
rect 6552 5034 6604 5040
rect 5448 5024 5500 5030
rect 5448 4966 5500 4972
rect 5460 4622 5488 4966
rect 5448 4616 5500 4622
rect 5448 4558 5500 4564
rect 6144 4380 6452 4400
rect 6144 4378 6150 4380
rect 6206 4378 6230 4380
rect 6286 4378 6310 4380
rect 6366 4378 6390 4380
rect 6446 4378 6452 4380
rect 6206 4326 6208 4378
rect 6388 4326 6390 4378
rect 6144 4324 6150 4326
rect 6206 4324 6230 4326
rect 6286 4324 6310 4326
rect 6366 4324 6390 4326
rect 6446 4324 6452 4326
rect 6144 4304 6452 4324
rect 5816 3936 5868 3942
rect 5816 3878 5868 3884
rect 5828 3534 5856 3878
rect 5816 3528 5868 3534
rect 5816 3470 5868 3476
rect 6144 3292 6452 3312
rect 6144 3290 6150 3292
rect 6206 3290 6230 3292
rect 6286 3290 6310 3292
rect 6366 3290 6390 3292
rect 6446 3290 6452 3292
rect 6206 3238 6208 3290
rect 6388 3238 6390 3290
rect 6144 3236 6150 3238
rect 6206 3236 6230 3238
rect 6286 3236 6310 3238
rect 6366 3236 6390 3238
rect 6446 3236 6452 3238
rect 6144 3216 6452 3236
rect 6564 3194 6592 5034
rect 7024 4146 7052 5578
rect 7443 4924 7751 4944
rect 7443 4922 7449 4924
rect 7505 4922 7529 4924
rect 7585 4922 7609 4924
rect 7665 4922 7689 4924
rect 7745 4922 7751 4924
rect 7505 4870 7507 4922
rect 7687 4870 7689 4922
rect 7443 4868 7449 4870
rect 7505 4868 7529 4870
rect 7585 4868 7609 4870
rect 7665 4868 7689 4870
rect 7745 4868 7751 4870
rect 7443 4848 7751 4868
rect 7012 4140 7064 4146
rect 7012 4082 7064 4088
rect 7104 3936 7156 3942
rect 7104 3878 7156 3884
rect 6552 3188 6604 3194
rect 6552 3130 6604 3136
rect 2136 2644 2188 2650
rect 2136 2586 2188 2592
rect 4252 2644 4304 2650
rect 4252 2586 4304 2592
rect 5264 2644 5316 2650
rect 5264 2586 5316 2592
rect 7116 2446 7144 3878
rect 7443 3836 7751 3856
rect 7443 3834 7449 3836
rect 7505 3834 7529 3836
rect 7585 3834 7609 3836
rect 7665 3834 7689 3836
rect 7745 3834 7751 3836
rect 7505 3782 7507 3834
rect 7687 3782 7689 3834
rect 7443 3780 7449 3782
rect 7505 3780 7529 3782
rect 7585 3780 7609 3782
rect 7665 3780 7689 3782
rect 7745 3780 7751 3782
rect 7443 3760 7751 3780
rect 8024 3392 8076 3398
rect 8024 3334 8076 3340
rect 8036 3097 8064 3334
rect 8022 3088 8078 3097
rect 8022 3023 8078 3032
rect 9588 3052 9640 3058
rect 9588 2994 9640 3000
rect 7443 2748 7751 2768
rect 7443 2746 7449 2748
rect 7505 2746 7529 2748
rect 7585 2746 7609 2748
rect 7665 2746 7689 2748
rect 7745 2746 7751 2748
rect 7505 2694 7507 2746
rect 7687 2694 7689 2746
rect 7443 2692 7449 2694
rect 7505 2692 7529 2694
rect 7585 2692 7609 2694
rect 7665 2692 7689 2694
rect 7745 2692 7751 2694
rect 7443 2672 7751 2692
rect 20 2440 72 2446
rect 20 2382 72 2388
rect 2412 2440 2464 2446
rect 2412 2382 2464 2388
rect 4804 2440 4856 2446
rect 4804 2382 4856 2388
rect 7104 2440 7156 2446
rect 7104 2382 7156 2388
rect 32 800 60 2382
rect 2424 800 2452 2382
rect 3547 2204 3855 2224
rect 3547 2202 3553 2204
rect 3609 2202 3633 2204
rect 3689 2202 3713 2204
rect 3769 2202 3793 2204
rect 3849 2202 3855 2204
rect 3609 2150 3611 2202
rect 3791 2150 3793 2202
rect 3547 2148 3553 2150
rect 3609 2148 3633 2150
rect 3689 2148 3713 2150
rect 3769 2148 3793 2150
rect 3849 2148 3855 2150
rect 3547 2128 3855 2148
rect 4816 800 4844 2382
rect 7196 2372 7248 2378
rect 7196 2314 7248 2320
rect 6144 2204 6452 2224
rect 6144 2202 6150 2204
rect 6206 2202 6230 2204
rect 6286 2202 6310 2204
rect 6366 2202 6390 2204
rect 6446 2202 6452 2204
rect 6206 2150 6208 2202
rect 6388 2150 6390 2202
rect 6144 2148 6150 2150
rect 6206 2148 6230 2150
rect 6286 2148 6310 2150
rect 6366 2148 6390 2150
rect 6446 2148 6452 2150
rect 6144 2128 6452 2148
rect 7208 800 7236 2314
rect 9600 800 9628 2994
rect 18 0 74 800
rect 2410 0 2466 800
rect 4802 0 4858 800
rect 7194 0 7250 800
rect 9586 0 9642 800
<< via2 >>
rect 2254 7098 2310 7100
rect 2334 7098 2390 7100
rect 2414 7098 2470 7100
rect 2494 7098 2550 7100
rect 2254 7046 2300 7098
rect 2300 7046 2310 7098
rect 2334 7046 2364 7098
rect 2364 7046 2376 7098
rect 2376 7046 2390 7098
rect 2414 7046 2428 7098
rect 2428 7046 2440 7098
rect 2440 7046 2470 7098
rect 2494 7046 2504 7098
rect 2504 7046 2550 7098
rect 2254 7044 2310 7046
rect 2334 7044 2390 7046
rect 2414 7044 2470 7046
rect 2494 7044 2550 7046
rect 1398 6840 1454 6896
rect 3553 7642 3609 7644
rect 3633 7642 3689 7644
rect 3713 7642 3769 7644
rect 3793 7642 3849 7644
rect 3553 7590 3599 7642
rect 3599 7590 3609 7642
rect 3633 7590 3663 7642
rect 3663 7590 3675 7642
rect 3675 7590 3689 7642
rect 3713 7590 3727 7642
rect 3727 7590 3739 7642
rect 3739 7590 3769 7642
rect 3793 7590 3803 7642
rect 3803 7590 3849 7642
rect 3553 7588 3609 7590
rect 3633 7588 3689 7590
rect 3713 7588 3769 7590
rect 3793 7588 3849 7590
rect 6150 7642 6206 7644
rect 6230 7642 6286 7644
rect 6310 7642 6366 7644
rect 6390 7642 6446 7644
rect 6150 7590 6196 7642
rect 6196 7590 6206 7642
rect 6230 7590 6260 7642
rect 6260 7590 6272 7642
rect 6272 7590 6286 7642
rect 6310 7590 6324 7642
rect 6324 7590 6336 7642
rect 6336 7590 6366 7642
rect 6390 7590 6400 7642
rect 6400 7590 6446 7642
rect 6150 7588 6206 7590
rect 6230 7588 6286 7590
rect 6310 7588 6366 7590
rect 6390 7588 6446 7590
rect 3553 6554 3609 6556
rect 3633 6554 3689 6556
rect 3713 6554 3769 6556
rect 3793 6554 3849 6556
rect 3553 6502 3599 6554
rect 3599 6502 3609 6554
rect 3633 6502 3663 6554
rect 3663 6502 3675 6554
rect 3675 6502 3689 6554
rect 3713 6502 3727 6554
rect 3727 6502 3739 6554
rect 3739 6502 3769 6554
rect 3793 6502 3803 6554
rect 3803 6502 3849 6554
rect 3553 6500 3609 6502
rect 3633 6500 3689 6502
rect 3713 6500 3769 6502
rect 3793 6500 3849 6502
rect 2254 6010 2310 6012
rect 2334 6010 2390 6012
rect 2414 6010 2470 6012
rect 2494 6010 2550 6012
rect 2254 5958 2300 6010
rect 2300 5958 2310 6010
rect 2334 5958 2364 6010
rect 2364 5958 2376 6010
rect 2376 5958 2390 6010
rect 2414 5958 2428 6010
rect 2428 5958 2440 6010
rect 2440 5958 2470 6010
rect 2494 5958 2504 6010
rect 2504 5958 2550 6010
rect 2254 5956 2310 5958
rect 2334 5956 2390 5958
rect 2414 5956 2470 5958
rect 2494 5956 2550 5958
rect 3553 5466 3609 5468
rect 3633 5466 3689 5468
rect 3713 5466 3769 5468
rect 3793 5466 3849 5468
rect 3553 5414 3599 5466
rect 3599 5414 3609 5466
rect 3633 5414 3663 5466
rect 3663 5414 3675 5466
rect 3675 5414 3689 5466
rect 3713 5414 3727 5466
rect 3727 5414 3739 5466
rect 3739 5414 3769 5466
rect 3793 5414 3803 5466
rect 3803 5414 3849 5466
rect 3553 5412 3609 5414
rect 3633 5412 3689 5414
rect 3713 5412 3769 5414
rect 3793 5412 3849 5414
rect 4852 7098 4908 7100
rect 4932 7098 4988 7100
rect 5012 7098 5068 7100
rect 5092 7098 5148 7100
rect 4852 7046 4898 7098
rect 4898 7046 4908 7098
rect 4932 7046 4962 7098
rect 4962 7046 4974 7098
rect 4974 7046 4988 7098
rect 5012 7046 5026 7098
rect 5026 7046 5038 7098
rect 5038 7046 5068 7098
rect 5092 7046 5102 7098
rect 5102 7046 5148 7098
rect 4852 7044 4908 7046
rect 4932 7044 4988 7046
rect 5012 7044 5068 7046
rect 5092 7044 5148 7046
rect 1398 3304 1454 3360
rect 2254 4922 2310 4924
rect 2334 4922 2390 4924
rect 2414 4922 2470 4924
rect 2494 4922 2550 4924
rect 2254 4870 2300 4922
rect 2300 4870 2310 4922
rect 2334 4870 2364 4922
rect 2364 4870 2376 4922
rect 2376 4870 2390 4922
rect 2414 4870 2428 4922
rect 2428 4870 2440 4922
rect 2440 4870 2470 4922
rect 2494 4870 2504 4922
rect 2504 4870 2550 4922
rect 2254 4868 2310 4870
rect 2334 4868 2390 4870
rect 2414 4868 2470 4870
rect 2494 4868 2550 4870
rect 4852 6010 4908 6012
rect 4932 6010 4988 6012
rect 5012 6010 5068 6012
rect 5092 6010 5148 6012
rect 4852 5958 4898 6010
rect 4898 5958 4908 6010
rect 4932 5958 4962 6010
rect 4962 5958 4974 6010
rect 4974 5958 4988 6010
rect 5012 5958 5026 6010
rect 5026 5958 5038 6010
rect 5038 5958 5068 6010
rect 5092 5958 5102 6010
rect 5102 5958 5148 6010
rect 4852 5956 4908 5958
rect 4932 5956 4988 5958
rect 5012 5956 5068 5958
rect 5092 5956 5148 5958
rect 4852 4922 4908 4924
rect 4932 4922 4988 4924
rect 5012 4922 5068 4924
rect 5092 4922 5148 4924
rect 4852 4870 4898 4922
rect 4898 4870 4908 4922
rect 4932 4870 4962 4922
rect 4962 4870 4974 4922
rect 4974 4870 4988 4922
rect 5012 4870 5026 4922
rect 5026 4870 5038 4922
rect 5038 4870 5068 4922
rect 5092 4870 5102 4922
rect 5102 4870 5148 4922
rect 4852 4868 4908 4870
rect 4932 4868 4988 4870
rect 5012 4868 5068 4870
rect 5092 4868 5148 4870
rect 6150 6554 6206 6556
rect 6230 6554 6286 6556
rect 6310 6554 6366 6556
rect 6390 6554 6446 6556
rect 6150 6502 6196 6554
rect 6196 6502 6206 6554
rect 6230 6502 6260 6554
rect 6260 6502 6272 6554
rect 6272 6502 6286 6554
rect 6310 6502 6324 6554
rect 6324 6502 6336 6554
rect 6336 6502 6366 6554
rect 6390 6502 6400 6554
rect 6400 6502 6446 6554
rect 6150 6500 6206 6502
rect 6230 6500 6286 6502
rect 6310 6500 6366 6502
rect 6390 6500 6446 6502
rect 7449 7098 7505 7100
rect 7529 7098 7585 7100
rect 7609 7098 7665 7100
rect 7689 7098 7745 7100
rect 7449 7046 7495 7098
rect 7495 7046 7505 7098
rect 7529 7046 7559 7098
rect 7559 7046 7571 7098
rect 7571 7046 7585 7098
rect 7609 7046 7623 7098
rect 7623 7046 7635 7098
rect 7635 7046 7665 7098
rect 7689 7046 7699 7098
rect 7699 7046 7745 7098
rect 7449 7044 7505 7046
rect 7529 7044 7585 7046
rect 7609 7044 7665 7046
rect 7689 7044 7745 7046
rect 7449 6010 7505 6012
rect 7529 6010 7585 6012
rect 7609 6010 7665 6012
rect 7689 6010 7745 6012
rect 7449 5958 7495 6010
rect 7495 5958 7505 6010
rect 7529 5958 7559 6010
rect 7559 5958 7571 6010
rect 7571 5958 7585 6010
rect 7609 5958 7623 6010
rect 7623 5958 7635 6010
rect 7635 5958 7665 6010
rect 7689 5958 7699 6010
rect 7699 5958 7745 6010
rect 7449 5956 7505 5958
rect 7529 5956 7585 5958
rect 7609 5956 7665 5958
rect 7689 5956 7745 5958
rect 8022 6604 8024 6624
rect 8024 6604 8076 6624
rect 8076 6604 8078 6624
rect 8022 6568 8078 6604
rect 6150 5466 6206 5468
rect 6230 5466 6286 5468
rect 6310 5466 6366 5468
rect 6390 5466 6446 5468
rect 6150 5414 6196 5466
rect 6196 5414 6206 5466
rect 6230 5414 6260 5466
rect 6260 5414 6272 5466
rect 6272 5414 6286 5466
rect 6310 5414 6324 5466
rect 6324 5414 6336 5466
rect 6336 5414 6366 5466
rect 6390 5414 6400 5466
rect 6400 5414 6446 5466
rect 6150 5412 6206 5414
rect 6230 5412 6286 5414
rect 6310 5412 6366 5414
rect 6390 5412 6446 5414
rect 3553 4378 3609 4380
rect 3633 4378 3689 4380
rect 3713 4378 3769 4380
rect 3793 4378 3849 4380
rect 3553 4326 3599 4378
rect 3599 4326 3609 4378
rect 3633 4326 3663 4378
rect 3663 4326 3675 4378
rect 3675 4326 3689 4378
rect 3713 4326 3727 4378
rect 3727 4326 3739 4378
rect 3739 4326 3769 4378
rect 3793 4326 3803 4378
rect 3803 4326 3849 4378
rect 3553 4324 3609 4326
rect 3633 4324 3689 4326
rect 3713 4324 3769 4326
rect 3793 4324 3849 4326
rect 2254 3834 2310 3836
rect 2334 3834 2390 3836
rect 2414 3834 2470 3836
rect 2494 3834 2550 3836
rect 2254 3782 2300 3834
rect 2300 3782 2310 3834
rect 2334 3782 2364 3834
rect 2364 3782 2376 3834
rect 2376 3782 2390 3834
rect 2414 3782 2428 3834
rect 2428 3782 2440 3834
rect 2440 3782 2470 3834
rect 2494 3782 2504 3834
rect 2504 3782 2550 3834
rect 2254 3780 2310 3782
rect 2334 3780 2390 3782
rect 2414 3780 2470 3782
rect 2494 3780 2550 3782
rect 3553 3290 3609 3292
rect 3633 3290 3689 3292
rect 3713 3290 3769 3292
rect 3793 3290 3849 3292
rect 3553 3238 3599 3290
rect 3599 3238 3609 3290
rect 3633 3238 3663 3290
rect 3663 3238 3675 3290
rect 3675 3238 3689 3290
rect 3713 3238 3727 3290
rect 3727 3238 3739 3290
rect 3739 3238 3769 3290
rect 3793 3238 3803 3290
rect 3803 3238 3849 3290
rect 3553 3236 3609 3238
rect 3633 3236 3689 3238
rect 3713 3236 3769 3238
rect 3793 3236 3849 3238
rect 2254 2746 2310 2748
rect 2334 2746 2390 2748
rect 2414 2746 2470 2748
rect 2494 2746 2550 2748
rect 2254 2694 2300 2746
rect 2300 2694 2310 2746
rect 2334 2694 2364 2746
rect 2364 2694 2376 2746
rect 2376 2694 2390 2746
rect 2414 2694 2428 2746
rect 2428 2694 2440 2746
rect 2440 2694 2470 2746
rect 2494 2694 2504 2746
rect 2504 2694 2550 2746
rect 2254 2692 2310 2694
rect 2334 2692 2390 2694
rect 2414 2692 2470 2694
rect 2494 2692 2550 2694
rect 4852 3834 4908 3836
rect 4932 3834 4988 3836
rect 5012 3834 5068 3836
rect 5092 3834 5148 3836
rect 4852 3782 4898 3834
rect 4898 3782 4908 3834
rect 4932 3782 4962 3834
rect 4962 3782 4974 3834
rect 4974 3782 4988 3834
rect 5012 3782 5026 3834
rect 5026 3782 5038 3834
rect 5038 3782 5068 3834
rect 5092 3782 5102 3834
rect 5102 3782 5148 3834
rect 4852 3780 4908 3782
rect 4932 3780 4988 3782
rect 5012 3780 5068 3782
rect 5092 3780 5148 3782
rect 4852 2746 4908 2748
rect 4932 2746 4988 2748
rect 5012 2746 5068 2748
rect 5092 2746 5148 2748
rect 4852 2694 4898 2746
rect 4898 2694 4908 2746
rect 4932 2694 4962 2746
rect 4962 2694 4974 2746
rect 4974 2694 4988 2746
rect 5012 2694 5026 2746
rect 5026 2694 5038 2746
rect 5038 2694 5068 2746
rect 5092 2694 5102 2746
rect 5102 2694 5148 2746
rect 4852 2692 4908 2694
rect 4932 2692 4988 2694
rect 5012 2692 5068 2694
rect 5092 2692 5148 2694
rect 6150 4378 6206 4380
rect 6230 4378 6286 4380
rect 6310 4378 6366 4380
rect 6390 4378 6446 4380
rect 6150 4326 6196 4378
rect 6196 4326 6206 4378
rect 6230 4326 6260 4378
rect 6260 4326 6272 4378
rect 6272 4326 6286 4378
rect 6310 4326 6324 4378
rect 6324 4326 6336 4378
rect 6336 4326 6366 4378
rect 6390 4326 6400 4378
rect 6400 4326 6446 4378
rect 6150 4324 6206 4326
rect 6230 4324 6286 4326
rect 6310 4324 6366 4326
rect 6390 4324 6446 4326
rect 6150 3290 6206 3292
rect 6230 3290 6286 3292
rect 6310 3290 6366 3292
rect 6390 3290 6446 3292
rect 6150 3238 6196 3290
rect 6196 3238 6206 3290
rect 6230 3238 6260 3290
rect 6260 3238 6272 3290
rect 6272 3238 6286 3290
rect 6310 3238 6324 3290
rect 6324 3238 6336 3290
rect 6336 3238 6366 3290
rect 6390 3238 6400 3290
rect 6400 3238 6446 3290
rect 6150 3236 6206 3238
rect 6230 3236 6286 3238
rect 6310 3236 6366 3238
rect 6390 3236 6446 3238
rect 7449 4922 7505 4924
rect 7529 4922 7585 4924
rect 7609 4922 7665 4924
rect 7689 4922 7745 4924
rect 7449 4870 7495 4922
rect 7495 4870 7505 4922
rect 7529 4870 7559 4922
rect 7559 4870 7571 4922
rect 7571 4870 7585 4922
rect 7609 4870 7623 4922
rect 7623 4870 7635 4922
rect 7635 4870 7665 4922
rect 7689 4870 7699 4922
rect 7699 4870 7745 4922
rect 7449 4868 7505 4870
rect 7529 4868 7585 4870
rect 7609 4868 7665 4870
rect 7689 4868 7745 4870
rect 7449 3834 7505 3836
rect 7529 3834 7585 3836
rect 7609 3834 7665 3836
rect 7689 3834 7745 3836
rect 7449 3782 7495 3834
rect 7495 3782 7505 3834
rect 7529 3782 7559 3834
rect 7559 3782 7571 3834
rect 7571 3782 7585 3834
rect 7609 3782 7623 3834
rect 7623 3782 7635 3834
rect 7635 3782 7665 3834
rect 7689 3782 7699 3834
rect 7699 3782 7745 3834
rect 7449 3780 7505 3782
rect 7529 3780 7585 3782
rect 7609 3780 7665 3782
rect 7689 3780 7745 3782
rect 8022 3032 8078 3088
rect 7449 2746 7505 2748
rect 7529 2746 7585 2748
rect 7609 2746 7665 2748
rect 7689 2746 7745 2748
rect 7449 2694 7495 2746
rect 7495 2694 7505 2746
rect 7529 2694 7559 2746
rect 7559 2694 7571 2746
rect 7571 2694 7585 2746
rect 7609 2694 7623 2746
rect 7623 2694 7635 2746
rect 7635 2694 7665 2746
rect 7689 2694 7699 2746
rect 7699 2694 7745 2746
rect 7449 2692 7505 2694
rect 7529 2692 7585 2694
rect 7609 2692 7665 2694
rect 7689 2692 7745 2694
rect 3553 2202 3609 2204
rect 3633 2202 3689 2204
rect 3713 2202 3769 2204
rect 3793 2202 3849 2204
rect 3553 2150 3599 2202
rect 3599 2150 3609 2202
rect 3633 2150 3663 2202
rect 3663 2150 3675 2202
rect 3675 2150 3689 2202
rect 3713 2150 3727 2202
rect 3727 2150 3739 2202
rect 3739 2150 3769 2202
rect 3793 2150 3803 2202
rect 3803 2150 3849 2202
rect 3553 2148 3609 2150
rect 3633 2148 3689 2150
rect 3713 2148 3769 2150
rect 3793 2148 3849 2150
rect 6150 2202 6206 2204
rect 6230 2202 6286 2204
rect 6310 2202 6366 2204
rect 6390 2202 6446 2204
rect 6150 2150 6196 2202
rect 6196 2150 6206 2202
rect 6230 2150 6260 2202
rect 6260 2150 6272 2202
rect 6272 2150 6286 2202
rect 6310 2150 6324 2202
rect 6324 2150 6336 2202
rect 6336 2150 6366 2202
rect 6390 2150 6400 2202
rect 6400 2150 6446 2202
rect 6150 2148 6206 2150
rect 6230 2148 6286 2150
rect 6310 2148 6366 2150
rect 6390 2148 6446 2150
<< metal3 >>
rect 3541 7648 3861 7649
rect 3541 7584 3549 7648
rect 3613 7584 3629 7648
rect 3693 7584 3709 7648
rect 3773 7584 3789 7648
rect 3853 7584 3861 7648
rect 3541 7583 3861 7584
rect 6138 7648 6458 7649
rect 6138 7584 6146 7648
rect 6210 7584 6226 7648
rect 6290 7584 6306 7648
rect 6370 7584 6386 7648
rect 6450 7584 6458 7648
rect 6138 7583 6458 7584
rect 2242 7104 2562 7105
rect 2242 7040 2250 7104
rect 2314 7040 2330 7104
rect 2394 7040 2410 7104
rect 2474 7040 2490 7104
rect 2554 7040 2562 7104
rect 2242 7039 2562 7040
rect 4840 7104 5160 7105
rect 4840 7040 4848 7104
rect 4912 7040 4928 7104
rect 4992 7040 5008 7104
rect 5072 7040 5088 7104
rect 5152 7040 5160 7104
rect 4840 7039 5160 7040
rect 7437 7104 7757 7105
rect 7437 7040 7445 7104
rect 7509 7040 7525 7104
rect 7589 7040 7605 7104
rect 7669 7040 7685 7104
rect 7749 7040 7757 7104
rect 7437 7039 7757 7040
rect 0 6898 800 6928
rect 1393 6898 1459 6901
rect 0 6896 1459 6898
rect 0 6840 1398 6896
rect 1454 6840 1459 6896
rect 0 6838 1459 6840
rect 0 6808 800 6838
rect 1393 6835 1459 6838
rect 8017 6626 8083 6629
rect 9200 6626 10000 6656
rect 8017 6624 10000 6626
rect 8017 6568 8022 6624
rect 8078 6568 10000 6624
rect 8017 6566 10000 6568
rect 8017 6563 8083 6566
rect 3541 6560 3861 6561
rect 3541 6496 3549 6560
rect 3613 6496 3629 6560
rect 3693 6496 3709 6560
rect 3773 6496 3789 6560
rect 3853 6496 3861 6560
rect 3541 6495 3861 6496
rect 6138 6560 6458 6561
rect 6138 6496 6146 6560
rect 6210 6496 6226 6560
rect 6290 6496 6306 6560
rect 6370 6496 6386 6560
rect 6450 6496 6458 6560
rect 9200 6536 10000 6566
rect 6138 6495 6458 6496
rect 2242 6016 2562 6017
rect 2242 5952 2250 6016
rect 2314 5952 2330 6016
rect 2394 5952 2410 6016
rect 2474 5952 2490 6016
rect 2554 5952 2562 6016
rect 2242 5951 2562 5952
rect 4840 6016 5160 6017
rect 4840 5952 4848 6016
rect 4912 5952 4928 6016
rect 4992 5952 5008 6016
rect 5072 5952 5088 6016
rect 5152 5952 5160 6016
rect 4840 5951 5160 5952
rect 7437 6016 7757 6017
rect 7437 5952 7445 6016
rect 7509 5952 7525 6016
rect 7589 5952 7605 6016
rect 7669 5952 7685 6016
rect 7749 5952 7757 6016
rect 7437 5951 7757 5952
rect 3541 5472 3861 5473
rect 3541 5408 3549 5472
rect 3613 5408 3629 5472
rect 3693 5408 3709 5472
rect 3773 5408 3789 5472
rect 3853 5408 3861 5472
rect 3541 5407 3861 5408
rect 6138 5472 6458 5473
rect 6138 5408 6146 5472
rect 6210 5408 6226 5472
rect 6290 5408 6306 5472
rect 6370 5408 6386 5472
rect 6450 5408 6458 5472
rect 6138 5407 6458 5408
rect 2242 4928 2562 4929
rect 2242 4864 2250 4928
rect 2314 4864 2330 4928
rect 2394 4864 2410 4928
rect 2474 4864 2490 4928
rect 2554 4864 2562 4928
rect 2242 4863 2562 4864
rect 4840 4928 5160 4929
rect 4840 4864 4848 4928
rect 4912 4864 4928 4928
rect 4992 4864 5008 4928
rect 5072 4864 5088 4928
rect 5152 4864 5160 4928
rect 4840 4863 5160 4864
rect 7437 4928 7757 4929
rect 7437 4864 7445 4928
rect 7509 4864 7525 4928
rect 7589 4864 7605 4928
rect 7669 4864 7685 4928
rect 7749 4864 7757 4928
rect 7437 4863 7757 4864
rect 3541 4384 3861 4385
rect 3541 4320 3549 4384
rect 3613 4320 3629 4384
rect 3693 4320 3709 4384
rect 3773 4320 3789 4384
rect 3853 4320 3861 4384
rect 3541 4319 3861 4320
rect 6138 4384 6458 4385
rect 6138 4320 6146 4384
rect 6210 4320 6226 4384
rect 6290 4320 6306 4384
rect 6370 4320 6386 4384
rect 6450 4320 6458 4384
rect 6138 4319 6458 4320
rect 2242 3840 2562 3841
rect 2242 3776 2250 3840
rect 2314 3776 2330 3840
rect 2394 3776 2410 3840
rect 2474 3776 2490 3840
rect 2554 3776 2562 3840
rect 2242 3775 2562 3776
rect 4840 3840 5160 3841
rect 4840 3776 4848 3840
rect 4912 3776 4928 3840
rect 4992 3776 5008 3840
rect 5072 3776 5088 3840
rect 5152 3776 5160 3840
rect 4840 3775 5160 3776
rect 7437 3840 7757 3841
rect 7437 3776 7445 3840
rect 7509 3776 7525 3840
rect 7589 3776 7605 3840
rect 7669 3776 7685 3840
rect 7749 3776 7757 3840
rect 7437 3775 7757 3776
rect 0 3362 800 3392
rect 1393 3362 1459 3365
rect 0 3360 1459 3362
rect 0 3304 1398 3360
rect 1454 3304 1459 3360
rect 0 3302 1459 3304
rect 0 3272 800 3302
rect 1393 3299 1459 3302
rect 3541 3296 3861 3297
rect 3541 3232 3549 3296
rect 3613 3232 3629 3296
rect 3693 3232 3709 3296
rect 3773 3232 3789 3296
rect 3853 3232 3861 3296
rect 3541 3231 3861 3232
rect 6138 3296 6458 3297
rect 6138 3232 6146 3296
rect 6210 3232 6226 3296
rect 6290 3232 6306 3296
rect 6370 3232 6386 3296
rect 6450 3232 6458 3296
rect 6138 3231 6458 3232
rect 8017 3090 8083 3093
rect 9200 3090 10000 3120
rect 8017 3088 10000 3090
rect 8017 3032 8022 3088
rect 8078 3032 10000 3088
rect 8017 3030 10000 3032
rect 8017 3027 8083 3030
rect 9200 3000 10000 3030
rect 2242 2752 2562 2753
rect 2242 2688 2250 2752
rect 2314 2688 2330 2752
rect 2394 2688 2410 2752
rect 2474 2688 2490 2752
rect 2554 2688 2562 2752
rect 2242 2687 2562 2688
rect 4840 2752 5160 2753
rect 4840 2688 4848 2752
rect 4912 2688 4928 2752
rect 4992 2688 5008 2752
rect 5072 2688 5088 2752
rect 5152 2688 5160 2752
rect 4840 2687 5160 2688
rect 7437 2752 7757 2753
rect 7437 2688 7445 2752
rect 7509 2688 7525 2752
rect 7589 2688 7605 2752
rect 7669 2688 7685 2752
rect 7749 2688 7757 2752
rect 7437 2687 7757 2688
rect 3541 2208 3861 2209
rect 3541 2144 3549 2208
rect 3613 2144 3629 2208
rect 3693 2144 3709 2208
rect 3773 2144 3789 2208
rect 3853 2144 3861 2208
rect 3541 2143 3861 2144
rect 6138 2208 6458 2209
rect 6138 2144 6146 2208
rect 6210 2144 6226 2208
rect 6290 2144 6306 2208
rect 6370 2144 6386 2208
rect 6450 2144 6458 2208
rect 6138 2143 6458 2144
<< via3 >>
rect 3549 7644 3613 7648
rect 3549 7588 3553 7644
rect 3553 7588 3609 7644
rect 3609 7588 3613 7644
rect 3549 7584 3613 7588
rect 3629 7644 3693 7648
rect 3629 7588 3633 7644
rect 3633 7588 3689 7644
rect 3689 7588 3693 7644
rect 3629 7584 3693 7588
rect 3709 7644 3773 7648
rect 3709 7588 3713 7644
rect 3713 7588 3769 7644
rect 3769 7588 3773 7644
rect 3709 7584 3773 7588
rect 3789 7644 3853 7648
rect 3789 7588 3793 7644
rect 3793 7588 3849 7644
rect 3849 7588 3853 7644
rect 3789 7584 3853 7588
rect 6146 7644 6210 7648
rect 6146 7588 6150 7644
rect 6150 7588 6206 7644
rect 6206 7588 6210 7644
rect 6146 7584 6210 7588
rect 6226 7644 6290 7648
rect 6226 7588 6230 7644
rect 6230 7588 6286 7644
rect 6286 7588 6290 7644
rect 6226 7584 6290 7588
rect 6306 7644 6370 7648
rect 6306 7588 6310 7644
rect 6310 7588 6366 7644
rect 6366 7588 6370 7644
rect 6306 7584 6370 7588
rect 6386 7644 6450 7648
rect 6386 7588 6390 7644
rect 6390 7588 6446 7644
rect 6446 7588 6450 7644
rect 6386 7584 6450 7588
rect 2250 7100 2314 7104
rect 2250 7044 2254 7100
rect 2254 7044 2310 7100
rect 2310 7044 2314 7100
rect 2250 7040 2314 7044
rect 2330 7100 2394 7104
rect 2330 7044 2334 7100
rect 2334 7044 2390 7100
rect 2390 7044 2394 7100
rect 2330 7040 2394 7044
rect 2410 7100 2474 7104
rect 2410 7044 2414 7100
rect 2414 7044 2470 7100
rect 2470 7044 2474 7100
rect 2410 7040 2474 7044
rect 2490 7100 2554 7104
rect 2490 7044 2494 7100
rect 2494 7044 2550 7100
rect 2550 7044 2554 7100
rect 2490 7040 2554 7044
rect 4848 7100 4912 7104
rect 4848 7044 4852 7100
rect 4852 7044 4908 7100
rect 4908 7044 4912 7100
rect 4848 7040 4912 7044
rect 4928 7100 4992 7104
rect 4928 7044 4932 7100
rect 4932 7044 4988 7100
rect 4988 7044 4992 7100
rect 4928 7040 4992 7044
rect 5008 7100 5072 7104
rect 5008 7044 5012 7100
rect 5012 7044 5068 7100
rect 5068 7044 5072 7100
rect 5008 7040 5072 7044
rect 5088 7100 5152 7104
rect 5088 7044 5092 7100
rect 5092 7044 5148 7100
rect 5148 7044 5152 7100
rect 5088 7040 5152 7044
rect 7445 7100 7509 7104
rect 7445 7044 7449 7100
rect 7449 7044 7505 7100
rect 7505 7044 7509 7100
rect 7445 7040 7509 7044
rect 7525 7100 7589 7104
rect 7525 7044 7529 7100
rect 7529 7044 7585 7100
rect 7585 7044 7589 7100
rect 7525 7040 7589 7044
rect 7605 7100 7669 7104
rect 7605 7044 7609 7100
rect 7609 7044 7665 7100
rect 7665 7044 7669 7100
rect 7605 7040 7669 7044
rect 7685 7100 7749 7104
rect 7685 7044 7689 7100
rect 7689 7044 7745 7100
rect 7745 7044 7749 7100
rect 7685 7040 7749 7044
rect 3549 6556 3613 6560
rect 3549 6500 3553 6556
rect 3553 6500 3609 6556
rect 3609 6500 3613 6556
rect 3549 6496 3613 6500
rect 3629 6556 3693 6560
rect 3629 6500 3633 6556
rect 3633 6500 3689 6556
rect 3689 6500 3693 6556
rect 3629 6496 3693 6500
rect 3709 6556 3773 6560
rect 3709 6500 3713 6556
rect 3713 6500 3769 6556
rect 3769 6500 3773 6556
rect 3709 6496 3773 6500
rect 3789 6556 3853 6560
rect 3789 6500 3793 6556
rect 3793 6500 3849 6556
rect 3849 6500 3853 6556
rect 3789 6496 3853 6500
rect 6146 6556 6210 6560
rect 6146 6500 6150 6556
rect 6150 6500 6206 6556
rect 6206 6500 6210 6556
rect 6146 6496 6210 6500
rect 6226 6556 6290 6560
rect 6226 6500 6230 6556
rect 6230 6500 6286 6556
rect 6286 6500 6290 6556
rect 6226 6496 6290 6500
rect 6306 6556 6370 6560
rect 6306 6500 6310 6556
rect 6310 6500 6366 6556
rect 6366 6500 6370 6556
rect 6306 6496 6370 6500
rect 6386 6556 6450 6560
rect 6386 6500 6390 6556
rect 6390 6500 6446 6556
rect 6446 6500 6450 6556
rect 6386 6496 6450 6500
rect 2250 6012 2314 6016
rect 2250 5956 2254 6012
rect 2254 5956 2310 6012
rect 2310 5956 2314 6012
rect 2250 5952 2314 5956
rect 2330 6012 2394 6016
rect 2330 5956 2334 6012
rect 2334 5956 2390 6012
rect 2390 5956 2394 6012
rect 2330 5952 2394 5956
rect 2410 6012 2474 6016
rect 2410 5956 2414 6012
rect 2414 5956 2470 6012
rect 2470 5956 2474 6012
rect 2410 5952 2474 5956
rect 2490 6012 2554 6016
rect 2490 5956 2494 6012
rect 2494 5956 2550 6012
rect 2550 5956 2554 6012
rect 2490 5952 2554 5956
rect 4848 6012 4912 6016
rect 4848 5956 4852 6012
rect 4852 5956 4908 6012
rect 4908 5956 4912 6012
rect 4848 5952 4912 5956
rect 4928 6012 4992 6016
rect 4928 5956 4932 6012
rect 4932 5956 4988 6012
rect 4988 5956 4992 6012
rect 4928 5952 4992 5956
rect 5008 6012 5072 6016
rect 5008 5956 5012 6012
rect 5012 5956 5068 6012
rect 5068 5956 5072 6012
rect 5008 5952 5072 5956
rect 5088 6012 5152 6016
rect 5088 5956 5092 6012
rect 5092 5956 5148 6012
rect 5148 5956 5152 6012
rect 5088 5952 5152 5956
rect 7445 6012 7509 6016
rect 7445 5956 7449 6012
rect 7449 5956 7505 6012
rect 7505 5956 7509 6012
rect 7445 5952 7509 5956
rect 7525 6012 7589 6016
rect 7525 5956 7529 6012
rect 7529 5956 7585 6012
rect 7585 5956 7589 6012
rect 7525 5952 7589 5956
rect 7605 6012 7669 6016
rect 7605 5956 7609 6012
rect 7609 5956 7665 6012
rect 7665 5956 7669 6012
rect 7605 5952 7669 5956
rect 7685 6012 7749 6016
rect 7685 5956 7689 6012
rect 7689 5956 7745 6012
rect 7745 5956 7749 6012
rect 7685 5952 7749 5956
rect 3549 5468 3613 5472
rect 3549 5412 3553 5468
rect 3553 5412 3609 5468
rect 3609 5412 3613 5468
rect 3549 5408 3613 5412
rect 3629 5468 3693 5472
rect 3629 5412 3633 5468
rect 3633 5412 3689 5468
rect 3689 5412 3693 5468
rect 3629 5408 3693 5412
rect 3709 5468 3773 5472
rect 3709 5412 3713 5468
rect 3713 5412 3769 5468
rect 3769 5412 3773 5468
rect 3709 5408 3773 5412
rect 3789 5468 3853 5472
rect 3789 5412 3793 5468
rect 3793 5412 3849 5468
rect 3849 5412 3853 5468
rect 3789 5408 3853 5412
rect 6146 5468 6210 5472
rect 6146 5412 6150 5468
rect 6150 5412 6206 5468
rect 6206 5412 6210 5468
rect 6146 5408 6210 5412
rect 6226 5468 6290 5472
rect 6226 5412 6230 5468
rect 6230 5412 6286 5468
rect 6286 5412 6290 5468
rect 6226 5408 6290 5412
rect 6306 5468 6370 5472
rect 6306 5412 6310 5468
rect 6310 5412 6366 5468
rect 6366 5412 6370 5468
rect 6306 5408 6370 5412
rect 6386 5468 6450 5472
rect 6386 5412 6390 5468
rect 6390 5412 6446 5468
rect 6446 5412 6450 5468
rect 6386 5408 6450 5412
rect 2250 4924 2314 4928
rect 2250 4868 2254 4924
rect 2254 4868 2310 4924
rect 2310 4868 2314 4924
rect 2250 4864 2314 4868
rect 2330 4924 2394 4928
rect 2330 4868 2334 4924
rect 2334 4868 2390 4924
rect 2390 4868 2394 4924
rect 2330 4864 2394 4868
rect 2410 4924 2474 4928
rect 2410 4868 2414 4924
rect 2414 4868 2470 4924
rect 2470 4868 2474 4924
rect 2410 4864 2474 4868
rect 2490 4924 2554 4928
rect 2490 4868 2494 4924
rect 2494 4868 2550 4924
rect 2550 4868 2554 4924
rect 2490 4864 2554 4868
rect 4848 4924 4912 4928
rect 4848 4868 4852 4924
rect 4852 4868 4908 4924
rect 4908 4868 4912 4924
rect 4848 4864 4912 4868
rect 4928 4924 4992 4928
rect 4928 4868 4932 4924
rect 4932 4868 4988 4924
rect 4988 4868 4992 4924
rect 4928 4864 4992 4868
rect 5008 4924 5072 4928
rect 5008 4868 5012 4924
rect 5012 4868 5068 4924
rect 5068 4868 5072 4924
rect 5008 4864 5072 4868
rect 5088 4924 5152 4928
rect 5088 4868 5092 4924
rect 5092 4868 5148 4924
rect 5148 4868 5152 4924
rect 5088 4864 5152 4868
rect 7445 4924 7509 4928
rect 7445 4868 7449 4924
rect 7449 4868 7505 4924
rect 7505 4868 7509 4924
rect 7445 4864 7509 4868
rect 7525 4924 7589 4928
rect 7525 4868 7529 4924
rect 7529 4868 7585 4924
rect 7585 4868 7589 4924
rect 7525 4864 7589 4868
rect 7605 4924 7669 4928
rect 7605 4868 7609 4924
rect 7609 4868 7665 4924
rect 7665 4868 7669 4924
rect 7605 4864 7669 4868
rect 7685 4924 7749 4928
rect 7685 4868 7689 4924
rect 7689 4868 7745 4924
rect 7745 4868 7749 4924
rect 7685 4864 7749 4868
rect 3549 4380 3613 4384
rect 3549 4324 3553 4380
rect 3553 4324 3609 4380
rect 3609 4324 3613 4380
rect 3549 4320 3613 4324
rect 3629 4380 3693 4384
rect 3629 4324 3633 4380
rect 3633 4324 3689 4380
rect 3689 4324 3693 4380
rect 3629 4320 3693 4324
rect 3709 4380 3773 4384
rect 3709 4324 3713 4380
rect 3713 4324 3769 4380
rect 3769 4324 3773 4380
rect 3709 4320 3773 4324
rect 3789 4380 3853 4384
rect 3789 4324 3793 4380
rect 3793 4324 3849 4380
rect 3849 4324 3853 4380
rect 3789 4320 3853 4324
rect 6146 4380 6210 4384
rect 6146 4324 6150 4380
rect 6150 4324 6206 4380
rect 6206 4324 6210 4380
rect 6146 4320 6210 4324
rect 6226 4380 6290 4384
rect 6226 4324 6230 4380
rect 6230 4324 6286 4380
rect 6286 4324 6290 4380
rect 6226 4320 6290 4324
rect 6306 4380 6370 4384
rect 6306 4324 6310 4380
rect 6310 4324 6366 4380
rect 6366 4324 6370 4380
rect 6306 4320 6370 4324
rect 6386 4380 6450 4384
rect 6386 4324 6390 4380
rect 6390 4324 6446 4380
rect 6446 4324 6450 4380
rect 6386 4320 6450 4324
rect 2250 3836 2314 3840
rect 2250 3780 2254 3836
rect 2254 3780 2310 3836
rect 2310 3780 2314 3836
rect 2250 3776 2314 3780
rect 2330 3836 2394 3840
rect 2330 3780 2334 3836
rect 2334 3780 2390 3836
rect 2390 3780 2394 3836
rect 2330 3776 2394 3780
rect 2410 3836 2474 3840
rect 2410 3780 2414 3836
rect 2414 3780 2470 3836
rect 2470 3780 2474 3836
rect 2410 3776 2474 3780
rect 2490 3836 2554 3840
rect 2490 3780 2494 3836
rect 2494 3780 2550 3836
rect 2550 3780 2554 3836
rect 2490 3776 2554 3780
rect 4848 3836 4912 3840
rect 4848 3780 4852 3836
rect 4852 3780 4908 3836
rect 4908 3780 4912 3836
rect 4848 3776 4912 3780
rect 4928 3836 4992 3840
rect 4928 3780 4932 3836
rect 4932 3780 4988 3836
rect 4988 3780 4992 3836
rect 4928 3776 4992 3780
rect 5008 3836 5072 3840
rect 5008 3780 5012 3836
rect 5012 3780 5068 3836
rect 5068 3780 5072 3836
rect 5008 3776 5072 3780
rect 5088 3836 5152 3840
rect 5088 3780 5092 3836
rect 5092 3780 5148 3836
rect 5148 3780 5152 3836
rect 5088 3776 5152 3780
rect 7445 3836 7509 3840
rect 7445 3780 7449 3836
rect 7449 3780 7505 3836
rect 7505 3780 7509 3836
rect 7445 3776 7509 3780
rect 7525 3836 7589 3840
rect 7525 3780 7529 3836
rect 7529 3780 7585 3836
rect 7585 3780 7589 3836
rect 7525 3776 7589 3780
rect 7605 3836 7669 3840
rect 7605 3780 7609 3836
rect 7609 3780 7665 3836
rect 7665 3780 7669 3836
rect 7605 3776 7669 3780
rect 7685 3836 7749 3840
rect 7685 3780 7689 3836
rect 7689 3780 7745 3836
rect 7745 3780 7749 3836
rect 7685 3776 7749 3780
rect 3549 3292 3613 3296
rect 3549 3236 3553 3292
rect 3553 3236 3609 3292
rect 3609 3236 3613 3292
rect 3549 3232 3613 3236
rect 3629 3292 3693 3296
rect 3629 3236 3633 3292
rect 3633 3236 3689 3292
rect 3689 3236 3693 3292
rect 3629 3232 3693 3236
rect 3709 3292 3773 3296
rect 3709 3236 3713 3292
rect 3713 3236 3769 3292
rect 3769 3236 3773 3292
rect 3709 3232 3773 3236
rect 3789 3292 3853 3296
rect 3789 3236 3793 3292
rect 3793 3236 3849 3292
rect 3849 3236 3853 3292
rect 3789 3232 3853 3236
rect 6146 3292 6210 3296
rect 6146 3236 6150 3292
rect 6150 3236 6206 3292
rect 6206 3236 6210 3292
rect 6146 3232 6210 3236
rect 6226 3292 6290 3296
rect 6226 3236 6230 3292
rect 6230 3236 6286 3292
rect 6286 3236 6290 3292
rect 6226 3232 6290 3236
rect 6306 3292 6370 3296
rect 6306 3236 6310 3292
rect 6310 3236 6366 3292
rect 6366 3236 6370 3292
rect 6306 3232 6370 3236
rect 6386 3292 6450 3296
rect 6386 3236 6390 3292
rect 6390 3236 6446 3292
rect 6446 3236 6450 3292
rect 6386 3232 6450 3236
rect 2250 2748 2314 2752
rect 2250 2692 2254 2748
rect 2254 2692 2310 2748
rect 2310 2692 2314 2748
rect 2250 2688 2314 2692
rect 2330 2748 2394 2752
rect 2330 2692 2334 2748
rect 2334 2692 2390 2748
rect 2390 2692 2394 2748
rect 2330 2688 2394 2692
rect 2410 2748 2474 2752
rect 2410 2692 2414 2748
rect 2414 2692 2470 2748
rect 2470 2692 2474 2748
rect 2410 2688 2474 2692
rect 2490 2748 2554 2752
rect 2490 2692 2494 2748
rect 2494 2692 2550 2748
rect 2550 2692 2554 2748
rect 2490 2688 2554 2692
rect 4848 2748 4912 2752
rect 4848 2692 4852 2748
rect 4852 2692 4908 2748
rect 4908 2692 4912 2748
rect 4848 2688 4912 2692
rect 4928 2748 4992 2752
rect 4928 2692 4932 2748
rect 4932 2692 4988 2748
rect 4988 2692 4992 2748
rect 4928 2688 4992 2692
rect 5008 2748 5072 2752
rect 5008 2692 5012 2748
rect 5012 2692 5068 2748
rect 5068 2692 5072 2748
rect 5008 2688 5072 2692
rect 5088 2748 5152 2752
rect 5088 2692 5092 2748
rect 5092 2692 5148 2748
rect 5148 2692 5152 2748
rect 5088 2688 5152 2692
rect 7445 2748 7509 2752
rect 7445 2692 7449 2748
rect 7449 2692 7505 2748
rect 7505 2692 7509 2748
rect 7445 2688 7509 2692
rect 7525 2748 7589 2752
rect 7525 2692 7529 2748
rect 7529 2692 7585 2748
rect 7585 2692 7589 2748
rect 7525 2688 7589 2692
rect 7605 2748 7669 2752
rect 7605 2692 7609 2748
rect 7609 2692 7665 2748
rect 7665 2692 7669 2748
rect 7605 2688 7669 2692
rect 7685 2748 7749 2752
rect 7685 2692 7689 2748
rect 7689 2692 7745 2748
rect 7745 2692 7749 2748
rect 7685 2688 7749 2692
rect 3549 2204 3613 2208
rect 3549 2148 3553 2204
rect 3553 2148 3609 2204
rect 3609 2148 3613 2204
rect 3549 2144 3613 2148
rect 3629 2204 3693 2208
rect 3629 2148 3633 2204
rect 3633 2148 3689 2204
rect 3689 2148 3693 2204
rect 3629 2144 3693 2148
rect 3709 2204 3773 2208
rect 3709 2148 3713 2204
rect 3713 2148 3769 2204
rect 3769 2148 3773 2204
rect 3709 2144 3773 2148
rect 3789 2204 3853 2208
rect 3789 2148 3793 2204
rect 3793 2148 3849 2204
rect 3849 2148 3853 2204
rect 3789 2144 3853 2148
rect 6146 2204 6210 2208
rect 6146 2148 6150 2204
rect 6150 2148 6206 2204
rect 6206 2148 6210 2204
rect 6146 2144 6210 2148
rect 6226 2204 6290 2208
rect 6226 2148 6230 2204
rect 6230 2148 6286 2204
rect 6286 2148 6290 2204
rect 6226 2144 6290 2148
rect 6306 2204 6370 2208
rect 6306 2148 6310 2204
rect 6310 2148 6366 2204
rect 6366 2148 6370 2204
rect 6306 2144 6370 2148
rect 6386 2204 6450 2208
rect 6386 2148 6390 2204
rect 6390 2148 6446 2204
rect 6446 2148 6450 2204
rect 6386 2144 6450 2148
<< metal4 >>
rect 2242 7104 2563 7664
rect 2242 7040 2250 7104
rect 2314 7040 2330 7104
rect 2394 7040 2410 7104
rect 2474 7040 2490 7104
rect 2554 7040 2563 7104
rect 2242 6952 2563 7040
rect 2242 6716 2284 6952
rect 2520 6716 2563 6952
rect 2242 6016 2563 6716
rect 2242 5952 2250 6016
rect 2314 5952 2330 6016
rect 2394 5952 2410 6016
rect 2474 5952 2490 6016
rect 2554 5952 2563 6016
rect 2242 5070 2563 5952
rect 2242 4928 2284 5070
rect 2520 4928 2563 5070
rect 2242 4864 2250 4928
rect 2554 4864 2563 4928
rect 2242 4834 2284 4864
rect 2520 4834 2563 4864
rect 2242 3840 2563 4834
rect 2242 3776 2250 3840
rect 2314 3776 2330 3840
rect 2394 3776 2410 3840
rect 2474 3776 2490 3840
rect 2554 3776 2563 3840
rect 2242 3187 2563 3776
rect 2242 2951 2284 3187
rect 2520 2951 2563 3187
rect 2242 2752 2563 2951
rect 2242 2688 2250 2752
rect 2314 2688 2330 2752
rect 2394 2688 2410 2752
rect 2474 2688 2490 2752
rect 2554 2688 2563 2752
rect 2242 2128 2563 2688
rect 3541 7648 3861 7664
rect 3541 7584 3549 7648
rect 3613 7584 3629 7648
rect 3693 7584 3709 7648
rect 3773 7584 3789 7648
rect 3853 7584 3861 7648
rect 3541 6560 3861 7584
rect 3541 6496 3549 6560
rect 3613 6496 3629 6560
rect 3693 6496 3709 6560
rect 3773 6496 3789 6560
rect 3853 6496 3861 6560
rect 3541 6011 3861 6496
rect 3541 5775 3583 6011
rect 3819 5775 3861 6011
rect 3541 5472 3861 5775
rect 3541 5408 3549 5472
rect 3613 5408 3629 5472
rect 3693 5408 3709 5472
rect 3773 5408 3789 5472
rect 3853 5408 3861 5472
rect 3541 4384 3861 5408
rect 3541 4320 3549 4384
rect 3613 4320 3629 4384
rect 3693 4320 3709 4384
rect 3773 4320 3789 4384
rect 3853 4320 3861 4384
rect 3541 4128 3861 4320
rect 3541 3892 3583 4128
rect 3819 3892 3861 4128
rect 3541 3296 3861 3892
rect 3541 3232 3549 3296
rect 3613 3232 3629 3296
rect 3693 3232 3709 3296
rect 3773 3232 3789 3296
rect 3853 3232 3861 3296
rect 3541 2208 3861 3232
rect 3541 2144 3549 2208
rect 3613 2144 3629 2208
rect 3693 2144 3709 2208
rect 3773 2144 3789 2208
rect 3853 2144 3861 2208
rect 3541 2128 3861 2144
rect 4840 7104 5160 7664
rect 4840 7040 4848 7104
rect 4912 7040 4928 7104
rect 4992 7040 5008 7104
rect 5072 7040 5088 7104
rect 5152 7040 5160 7104
rect 4840 6952 5160 7040
rect 4840 6716 4882 6952
rect 5118 6716 5160 6952
rect 4840 6016 5160 6716
rect 4840 5952 4848 6016
rect 4912 5952 4928 6016
rect 4992 5952 5008 6016
rect 5072 5952 5088 6016
rect 5152 5952 5160 6016
rect 4840 5070 5160 5952
rect 4840 4928 4882 5070
rect 5118 4928 5160 5070
rect 4840 4864 4848 4928
rect 5152 4864 5160 4928
rect 4840 4834 4882 4864
rect 5118 4834 5160 4864
rect 4840 3840 5160 4834
rect 4840 3776 4848 3840
rect 4912 3776 4928 3840
rect 4992 3776 5008 3840
rect 5072 3776 5088 3840
rect 5152 3776 5160 3840
rect 4840 3187 5160 3776
rect 4840 2951 4882 3187
rect 5118 2951 5160 3187
rect 4840 2752 5160 2951
rect 4840 2688 4848 2752
rect 4912 2688 4928 2752
rect 4992 2688 5008 2752
rect 5072 2688 5088 2752
rect 5152 2688 5160 2752
rect 4840 2128 5160 2688
rect 6138 7648 6458 7664
rect 6138 7584 6146 7648
rect 6210 7584 6226 7648
rect 6290 7584 6306 7648
rect 6370 7584 6386 7648
rect 6450 7584 6458 7648
rect 6138 6560 6458 7584
rect 6138 6496 6146 6560
rect 6210 6496 6226 6560
rect 6290 6496 6306 6560
rect 6370 6496 6386 6560
rect 6450 6496 6458 6560
rect 6138 6011 6458 6496
rect 6138 5775 6180 6011
rect 6416 5775 6458 6011
rect 6138 5472 6458 5775
rect 6138 5408 6146 5472
rect 6210 5408 6226 5472
rect 6290 5408 6306 5472
rect 6370 5408 6386 5472
rect 6450 5408 6458 5472
rect 6138 4384 6458 5408
rect 6138 4320 6146 4384
rect 6210 4320 6226 4384
rect 6290 4320 6306 4384
rect 6370 4320 6386 4384
rect 6450 4320 6458 4384
rect 6138 4128 6458 4320
rect 6138 3892 6180 4128
rect 6416 3892 6458 4128
rect 6138 3296 6458 3892
rect 6138 3232 6146 3296
rect 6210 3232 6226 3296
rect 6290 3232 6306 3296
rect 6370 3232 6386 3296
rect 6450 3232 6458 3296
rect 6138 2208 6458 3232
rect 6138 2144 6146 2208
rect 6210 2144 6226 2208
rect 6290 2144 6306 2208
rect 6370 2144 6386 2208
rect 6450 2144 6458 2208
rect 6138 2128 6458 2144
rect 7437 7104 7757 7664
rect 7437 7040 7445 7104
rect 7509 7040 7525 7104
rect 7589 7040 7605 7104
rect 7669 7040 7685 7104
rect 7749 7040 7757 7104
rect 7437 6952 7757 7040
rect 7437 6716 7479 6952
rect 7715 6716 7757 6952
rect 7437 6016 7757 6716
rect 7437 5952 7445 6016
rect 7509 5952 7525 6016
rect 7589 5952 7605 6016
rect 7669 5952 7685 6016
rect 7749 5952 7757 6016
rect 7437 5070 7757 5952
rect 7437 4928 7479 5070
rect 7715 4928 7757 5070
rect 7437 4864 7445 4928
rect 7749 4864 7757 4928
rect 7437 4834 7479 4864
rect 7715 4834 7757 4864
rect 7437 3840 7757 4834
rect 7437 3776 7445 3840
rect 7509 3776 7525 3840
rect 7589 3776 7605 3840
rect 7669 3776 7685 3840
rect 7749 3776 7757 3840
rect 7437 3187 7757 3776
rect 7437 2951 7479 3187
rect 7715 2951 7757 3187
rect 7437 2752 7757 2951
rect 7437 2688 7445 2752
rect 7509 2688 7525 2752
rect 7589 2688 7605 2752
rect 7669 2688 7685 2752
rect 7749 2688 7757 2752
rect 7437 2128 7757 2688
<< via4 >>
rect 2284 6716 2520 6952
rect 2284 4928 2520 5070
rect 2284 4864 2314 4928
rect 2314 4864 2330 4928
rect 2330 4864 2394 4928
rect 2394 4864 2410 4928
rect 2410 4864 2474 4928
rect 2474 4864 2490 4928
rect 2490 4864 2520 4928
rect 2284 4834 2520 4864
rect 2284 2951 2520 3187
rect 3583 5775 3819 6011
rect 3583 3892 3819 4128
rect 4882 6716 5118 6952
rect 4882 4928 5118 5070
rect 4882 4864 4912 4928
rect 4912 4864 4928 4928
rect 4928 4864 4992 4928
rect 4992 4864 5008 4928
rect 5008 4864 5072 4928
rect 5072 4864 5088 4928
rect 5088 4864 5118 4928
rect 4882 4834 5118 4864
rect 4882 2951 5118 3187
rect 6180 5775 6416 6011
rect 6180 3892 6416 4128
rect 7479 6716 7715 6952
rect 7479 4928 7715 5070
rect 7479 4864 7509 4928
rect 7509 4864 7525 4928
rect 7525 4864 7589 4928
rect 7589 4864 7605 4928
rect 7605 4864 7669 4928
rect 7669 4864 7685 4928
rect 7685 4864 7715 4928
rect 7479 4834 7715 4864
rect 7479 2951 7715 3187
<< metal5 >>
rect 1104 6952 8832 6994
rect 1104 6716 2284 6952
rect 2520 6716 4882 6952
rect 5118 6716 7479 6952
rect 7715 6716 8832 6952
rect 1104 6674 8832 6716
rect 1104 6011 8832 6053
rect 1104 5775 3583 6011
rect 3819 5775 6180 6011
rect 6416 5775 8832 6011
rect 1104 5733 8832 5775
rect 1104 5070 8832 5112
rect 1104 4834 2284 5070
rect 2520 4834 4882 5070
rect 5118 4834 7479 5070
rect 7715 4834 8832 5070
rect 1104 4792 8832 4834
rect 1104 4128 8832 4170
rect 1104 3892 3583 4128
rect 3819 3892 6180 4128
rect 6416 3892 8832 4128
rect 1104 3850 8832 3892
rect 1104 3187 8832 3229
rect 1104 2951 2284 3187
rect 2520 2951 4882 3187
rect 5118 2951 7479 3187
rect 7715 2951 8832 3187
rect 1104 2909 8832 2951
use sky130_fd_sc_hd__decap_8  FILLER_0_6 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1633346062
transform 1 0 1656 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_1_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1633346062
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1633346062
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1633346062
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input4 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1633346062
transform 1 0 1380 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1633346062
transform 1 0 2392 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18
timestamp 1633346062
transform 1 0 2760 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_1_15
timestamp 1633346062
transform 1 0 2484 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  input1
timestamp 1633346062
transform 1 0 2484 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1633346062
transform 1 0 3496 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_0_29
timestamp 1633346062
transform 1 0 3772 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_27
timestamp 1633346062
transform 1 0 3588 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_20 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1633346062
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_44
timestamp 1633346062
transform 1 0 5152 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_39
timestamp 1633346062
transform 1 0 4692 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_51 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1633346062
transform 1 0 5796 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input9
timestamp 1633346062
transform 1 0 4876 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_57
timestamp 1633346062
transform 1 0 6348 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_55
timestamp 1633346062
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_57
timestamp 1633346062
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_21
timestamp 1633346062
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_22
timestamp 1633346062
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_65
timestamp 1633346062
transform 1 0 7084 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_71
timestamp 1633346062
transform 1 0 7636 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_1_69
timestamp 1633346062
transform 1 0 7452 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_73
timestamp 1633346062
transform 1 0 7820 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_77
timestamp 1633346062
transform 1 0 8188 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input6
timestamp 1633346062
transform -1 0 8188 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output11 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1633346062
transform -1 0 7636 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_79
timestamp 1633346062
transform 1 0 8372 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1633346062
transform -1 0 8832 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1633346062
transform -1 0 8832 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_2_6
timestamp 1633346062
transform 1 0 1656 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1633346062
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input2 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1633346062
transform -1 0 1656 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_2_18
timestamp 1633346062
transform 1 0 2760 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_26
timestamp 1633346062
transform 1 0 3496 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_2_29
timestamp 1633346062
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_23
timestamp 1633346062
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_41
timestamp 1633346062
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_53
timestamp 1633346062
transform 1 0 5980 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_65
timestamp 1633346062
transform 1 0 7084 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_2_77
timestamp 1633346062
transform 1 0 8188 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output14
timestamp 1633346062
transform 1 0 7820 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1633346062
transform -1 0 8832 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_3_3
timestamp 1633346062
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1633346062
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_3_15
timestamp 1633346062
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_27
timestamp 1633346062
transform 1 0 3588 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_3_39
timestamp 1633346062
transform 1 0 4692 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__dlxtp_1  _30_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1633346062
transform 1 0 4784 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_52
timestamp 1633346062
transform 1 0 5888 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_57 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1633346062
transform 1 0 6348 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_63
timestamp 1633346062
transform 1 0 6900 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_24
timestamp 1633346062
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _27_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1633346062
transform 1 0 6992 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_3_67
timestamp 1633346062
transform 1 0 7268 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_3_79
timestamp 1633346062
transform 1 0 8372 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1633346062
transform -1 0 8832 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_4_3
timestamp 1633346062
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1633346062
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_4_15
timestamp 1633346062
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp 1633346062
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_29
timestamp 1633346062
transform 1 0 3772 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_33
timestamp 1633346062
transform 1 0 4140 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_37
timestamp 1633346062
transform 1 0 4508 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_25
timestamp 1633346062
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _25_
timestamp 1633346062
transform 1 0 4232 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_4_48
timestamp 1633346062
transform 1 0 5520 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  _15_
timestamp 1633346062
transform 1 0 5244 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_4_60
timestamp 1633346062
transform 1 0 6624 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_72
timestamp 1633346062
transform 1 0 7728 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_80
timestamp 1633346062
transform 1 0 8464 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1633346062
transform -1 0 8832 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_5_11
timestamp 1633346062
transform 1 0 2116 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_3
timestamp 1633346062
transform 1 0 1380 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1633346062
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _24_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1633346062
transform -1 0 2852 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__decap_6  FILLER_5_19
timestamp 1633346062
transform 1 0 2852 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _21_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1633346062
transform 1 0 3404 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__decap_6  FILLER_5_30
timestamp 1633346062
transform 1 0 3864 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _18_
timestamp 1633346062
transform -1 0 4692 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_5_39
timestamp 1633346062
transform 1 0 4692 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_5_51
timestamp 1633346062
transform 1 0 5796 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__or4_1  _14_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1633346062
transform 1 0 5244 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_55
timestamp 1633346062
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_60
timestamp 1633346062
transform 1 0 6624 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_26
timestamp 1633346062
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _20_
timestamp 1633346062
transform -1 0 6624 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_5_72
timestamp 1633346062
transform 1 0 7728 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_80
timestamp 1633346062
transform 1 0 8464 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1633346062
transform -1 0 8832 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_6_3
timestamp 1633346062
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_3
timestamp 1633346062
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1633346062
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1633346062
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_6_15
timestamp 1633346062
transform 1 0 2484 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_19
timestamp 1633346062
transform 1 0 2852 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_23
timestamp 1633346062
transform 1 0 3220 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_15
timestamp 1633346062
transform 1 0 2484 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_19
timestamp 1633346062
transform 1 0 2852 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_7_24
timestamp 1633346062
transform 1 0 3312 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _16_
timestamp 1633346062
transform 1 0 2944 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _17_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1633346062
transform -1 0 3312 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp 1633346062
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_6_29
timestamp 1633346062
transform 1 0 3772 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_27
timestamp 1633346062
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__a311o_1  _22_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1633346062
transform 1 0 4048 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__a41o_1  _26_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1633346062
transform -1 0 5060 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_6_43
timestamp 1633346062
transform 1 0 5060 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_6_50
timestamp 1633346062
transform 1 0 5704 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_40
timestamp 1633346062
transform 1 0 4784 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__nor2_1  _23_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1633346062
transform -1 0 5704 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_6_62
timestamp 1633346062
transform 1 0 6808 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_52
timestamp 1633346062
transform 1 0 5888 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_7_57
timestamp 1633346062
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_28
timestamp 1633346062
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_6_74
timestamp 1633346062
transform 1 0 7912 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_7_69
timestamp 1633346062
transform 1 0 7452 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_80
timestamp 1633346062
transform 1 0 8464 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1633346062
transform -1 0 8832 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1633346062
transform -1 0 8832 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_8_6
timestamp 1633346062
transform 1 0 1656 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1633346062
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1633346062
transform -1 0 1656 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_14
timestamp 1633346062
transform 1 0 2392 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_8_21
timestamp 1633346062
transform 1 0 3036 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  output13
timestamp 1633346062
transform -1 0 3036 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_27
timestamp 1633346062
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_8_29
timestamp 1633346062
transform 1 0 3772 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_37
timestamp 1633346062
transform 1 0 4508 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_29
timestamp 1633346062
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__o221ai_1  _19_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1633346062
transform 1 0 3864 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_8_44
timestamp 1633346062
transform 1 0 5152 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _13_
timestamp 1633346062
transform -1 0 5152 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_8_56
timestamp 1633346062
transform 1 0 6256 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_68
timestamp 1633346062
transform 1 0 7360 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_72
timestamp 1633346062
transform 1 0 7728 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_77
timestamp 1633346062
transform 1 0 8188 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output10
timestamp 1633346062
transform 1 0 7820 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1633346062
transform -1 0 8832 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_9_7
timestamp 1633346062
transform 1 0 1748 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1633346062
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__dlxtp_1  _28_
timestamp 1633346062
transform -1 0 3220 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_2  output12
timestamp 1633346062
transform -1 0 1748 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_23
timestamp 1633346062
transform 1 0 3220 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_27
timestamp 1633346062
transform 1 0 3588 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_30
timestamp 1633346062
transform 1 0 3680 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__dlxtp_1  _29_
timestamp 1633346062
transform -1 0 4876 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_41
timestamp 1633346062
transform 1 0 4876 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_9_48
timestamp 1633346062
transform 1 0 5520 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  input7
timestamp 1633346062
transform 1 0 5244 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_9_57
timestamp 1633346062
transform 1 0 6348 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_61
timestamp 1633346062
transform 1 0 6716 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_31
timestamp 1633346062
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input8
timestamp 1633346062
transform -1 0 7084 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_9_65
timestamp 1633346062
transform 1 0 7084 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_9_72
timestamp 1633346062
transform 1 0 7728 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  input5
timestamp 1633346062
transform -1 0 7728 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_9_80
timestamp 1633346062
transform 1 0 8464 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1633346062
transform -1 0 8832 0 -1 7616
box -38 -48 314 592
<< labels >>
rlabel metal5 s 1104 3850 8832 4170 6 VGND
port 0 nsew ground input
rlabel metal5 s 1104 5733 8832 6053 6 VGND
port 0 nsew ground input
rlabel metal4 s 3541 2128 3861 7664 6 VGND
port 0 nsew ground input
rlabel metal4 s 6138 2128 6458 7664 6 VGND
port 0 nsew ground input
rlabel metal5 s 1104 2909 8832 3229 6 VPWR
port 1 nsew power input
rlabel metal5 s 1104 4792 8832 5112 6 VPWR
port 1 nsew power input
rlabel metal5 s 1104 6674 8832 6994 6 VPWR
port 1 nsew power input
rlabel metal4 s 2243 2128 2563 7664 6 VPWR
port 1 nsew power input
rlabel metal4 s 4840 2128 5160 7664 6 VPWR
port 1 nsew power input
rlabel metal4 s 7437 2128 7757 7664 6 VPWR
port 1 nsew power input
rlabel metal2 s 2410 0 2466 800 6 en
port 2 nsew signal input
rlabel metal3 s 9200 6536 10000 6656 6 eno
port 3 nsew signal tristate
rlabel metal2 s 7194 0 7250 800 6 gs
port 4 nsew signal tristate
rlabel metal3 s 0 3272 800 3392 6 in[0]
port 5 nsew signal input
rlabel metal3 s 0 6808 800 6928 6 in[1]
port 6 nsew signal input
rlabel metal2 s 18 0 74 800 6 in[2]
port 7 nsew signal input
rlabel metal2 s 7378 9200 7434 10000 6 in[3]
port 8 nsew signal input
rlabel metal2 s 9586 0 9642 800 6 in[4]
port 9 nsew signal input
rlabel metal2 s 4986 9200 5042 10000 6 in[5]
port 10 nsew signal input
rlabel metal2 s 9770 9200 9826 10000 6 in[6]
port 11 nsew signal input
rlabel metal2 s 4802 0 4858 800 6 in[7]
port 12 nsew signal input
rlabel metal2 s 202 9200 258 10000 6 out[0]
port 13 nsew signal tristate
rlabel metal2 s 2594 9200 2650 10000 6 out[1]
port 14 nsew signal tristate
rlabel metal3 s 9200 3000 10000 3120 6 out[2]
port 15 nsew signal tristate
<< properties >>
string FIXED_BBOX 0 0 10000 10000
<< end >>
