magic
tech sky130A
magscale 1 2
timestamp 1634271525
<< obsli1 >>
rect 1104 2159 8832 7633
<< obsm1 >>
rect 14 2128 9830 7664
<< metal2 >>
rect 202 9200 258 10000
rect 2594 9200 2650 10000
rect 4986 9200 5042 10000
rect 7378 9200 7434 10000
rect 9770 9200 9826 10000
rect 18 0 74 800
rect 2410 0 2466 800
rect 4802 0 4858 800
rect 7194 0 7250 800
rect 9586 0 9642 800
<< obsm2 >>
rect 20 9144 146 9200
rect 314 9144 2538 9200
rect 2706 9144 4930 9200
rect 5098 9144 7322 9200
rect 7490 9144 9714 9200
rect 20 856 9824 9144
rect 130 800 2354 856
rect 2522 800 4746 856
rect 4914 800 7138 856
rect 7306 800 9530 856
rect 9698 800 9824 856
<< metal3 >>
rect 0 6808 800 6928
rect 9200 6536 10000 6656
rect 0 3272 800 3392
rect 9200 3000 10000 3120
<< obsm3 >>
rect 800 7008 9200 7649
rect 880 6736 9200 7008
rect 880 6728 9120 6736
rect 800 6456 9120 6728
rect 800 3472 9200 6456
rect 880 3200 9200 3472
rect 880 3192 9120 3200
rect 800 2920 9120 3192
rect 800 2143 9200 2920
<< metal4 >>
rect 2243 2128 2563 7664
rect 3541 2128 3861 7664
rect 4840 2128 5160 7664
rect 6138 2128 6458 7664
rect 7437 2128 7757 7664
<< metal5 >>
rect 1104 6674 8832 6994
rect 1104 5733 8832 6053
rect 1104 4792 8832 5112
rect 1104 3850 8832 4170
rect 1104 2909 8832 3229
<< labels >>
rlabel metal5 s 1104 3850 8832 4170 6 VGND
port 1 nsew ground input
rlabel metal5 s 1104 5733 8832 6053 6 VGND
port 1 nsew ground input
rlabel metal4 s 3541 2128 3861 7664 6 VGND
port 1 nsew ground input
rlabel metal4 s 6138 2128 6458 7664 6 VGND
port 1 nsew ground input
rlabel metal5 s 1104 2909 8832 3229 6 VPWR
port 2 nsew power input
rlabel metal5 s 1104 4792 8832 5112 6 VPWR
port 2 nsew power input
rlabel metal5 s 1104 6674 8832 6994 6 VPWR
port 2 nsew power input
rlabel metal4 s 2243 2128 2563 7664 6 VPWR
port 2 nsew power input
rlabel metal4 s 4840 2128 5160 7664 6 VPWR
port 2 nsew power input
rlabel metal4 s 7437 2128 7757 7664 6 VPWR
port 2 nsew power input
rlabel metal2 s 2410 0 2466 800 6 en
port 3 nsew signal input
rlabel metal3 s 9200 6536 10000 6656 6 eno
port 4 nsew signal output
rlabel metal2 s 7194 0 7250 800 6 gs
port 5 nsew signal output
rlabel metal3 s 0 3272 800 3392 6 in[0]
port 6 nsew signal input
rlabel metal3 s 0 6808 800 6928 6 in[1]
port 7 nsew signal input
rlabel metal2 s 18 0 74 800 6 in[2]
port 8 nsew signal input
rlabel metal2 s 7378 9200 7434 10000 6 in[3]
port 9 nsew signal input
rlabel metal2 s 9586 0 9642 800 6 in[4]
port 10 nsew signal input
rlabel metal2 s 4986 9200 5042 10000 6 in[5]
port 11 nsew signal input
rlabel metal2 s 9770 9200 9826 10000 6 in[6]
port 12 nsew signal input
rlabel metal2 s 4802 0 4858 800 6 in[7]
port 13 nsew signal input
rlabel metal2 s 202 9200 258 10000 6 out[0]
port 14 nsew signal output
rlabel metal2 s 2594 9200 2650 10000 6 out[1]
port 15 nsew signal output
rlabel metal3 s 9200 3000 10000 3120 6 out[2]
port 16 nsew signal output
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 10000 10000
string LEFview TRUE
string GDS_FILE /openLANE_flow/designs/dvsd_pe/runs/15-10_04-15/results/magic/dvsd_pe.gds
string GDS_END 190246
string GDS_START 93176
<< end >>

