magic
tech sky130A
magscale 1 2
timestamp 1633167455
<< obsli1 >>
rect 1104 2159 178848 117521
<< obsm1 >>
rect 14 2128 179846 117552
<< metal2 >>
rect 30746 119200 30802 120000
rect 67914 119200 67970 120000
rect 105266 119200 105322 120000
rect 142618 119200 142674 120000
rect 179786 119200 179842 120000
rect 18 0 74 800
rect 37186 0 37242 800
rect 74538 0 74594 800
rect 111890 0 111946 800
rect 149058 0 149114 800
<< obsm2 >>
rect 20 119144 30690 119200
rect 30858 119144 67858 119200
rect 68026 119144 105210 119200
rect 105378 119144 142562 119200
rect 142730 119144 179730 119200
rect 20 856 179840 119144
rect 130 800 37130 856
rect 37298 800 74482 856
rect 74650 800 111834 856
rect 112002 800 149002 856
rect 149170 800 179840 856
<< metal3 >>
rect 0 110168 800 110288
rect 179200 64744 180000 64864
rect 0 54952 800 55072
rect 179200 9528 180000 9648
<< obsm3 >>
rect 800 110368 179200 117537
rect 880 110088 179200 110368
rect 800 64944 179200 110088
rect 800 64664 179120 64944
rect 800 55152 179200 64664
rect 880 54872 179200 55152
rect 800 9728 179200 54872
rect 800 9448 179120 9728
rect 800 2143 179200 9448
<< metal4 >>
rect 4208 2128 4528 117552
rect 19568 2128 19888 117552
rect 34928 2128 35248 117552
rect 50288 2128 50608 117552
rect 65648 2128 65968 117552
rect 81008 2128 81328 117552
rect 96368 2128 96688 117552
rect 111728 2128 112048 117552
rect 127088 2128 127408 117552
rect 142448 2128 142768 117552
rect 157808 2128 158128 117552
rect 173168 2128 173488 117552
<< labels >>
rlabel metal4 s 19568 2128 19888 117552 6 VGND
port 1 nsew ground input
rlabel metal4 s 50288 2128 50608 117552 6 VGND
port 1 nsew ground input
rlabel metal4 s 81008 2128 81328 117552 6 VGND
port 1 nsew ground input
rlabel metal4 s 111728 2128 112048 117552 6 VGND
port 1 nsew ground input
rlabel metal4 s 142448 2128 142768 117552 6 VGND
port 1 nsew ground input
rlabel metal4 s 173168 2128 173488 117552 6 VGND
port 1 nsew ground input
rlabel metal4 s 4208 2128 4528 117552 6 VPWR
port 2 nsew power input
rlabel metal4 s 34928 2128 35248 117552 6 VPWR
port 2 nsew power input
rlabel metal4 s 65648 2128 65968 117552 6 VPWR
port 2 nsew power input
rlabel metal4 s 96368 2128 96688 117552 6 VPWR
port 2 nsew power input
rlabel metal4 s 127088 2128 127408 117552 6 VPWR
port 2 nsew power input
rlabel metal4 s 157808 2128 158128 117552 6 VPWR
port 2 nsew power input
rlabel metal2 s 37186 0 37242 800 6 io_en
port 3 nsew signal input
rlabel metal3 s 179200 64744 180000 64864 6 io_in[0]
port 4 nsew signal input
rlabel metal2 s 111890 0 111946 800 6 io_in[1]
port 5 nsew signal input
rlabel metal3 s 0 54952 800 55072 6 io_in[2]
port 6 nsew signal input
rlabel metal3 s 0 110168 800 110288 6 io_in[3]
port 7 nsew signal input
rlabel metal2 s 18 0 74 800 6 io_in[4]
port 8 nsew signal input
rlabel metal2 s 142618 119200 142674 120000 6 io_in[5]
port 9 nsew signal input
rlabel metal2 s 149058 0 149114 800 6 io_in[6]
port 10 nsew signal input
rlabel metal2 s 105266 119200 105322 120000 6 io_in[7]
port 11 nsew signal input
rlabel metal2 s 179786 119200 179842 120000 6 io_out[0]
port 12 nsew signal output
rlabel metal2 s 74538 0 74594 800 6 io_out[1]
port 13 nsew signal output
rlabel metal2 s 30746 119200 30802 120000 6 io_out[2]
port 14 nsew signal output
rlabel metal2 s 67914 119200 67970 120000 6 wb_eno
port 15 nsew signal output
rlabel metal3 s 179200 9528 180000 9648 6 wb_gs
port 16 nsew signal output
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 180000 120000
string LEFview TRUE
string GDS_FILE /project/openlane/user_proj_example/runs/user_proj_example/results/magic/user_proj_example.gds
string GDS_END 5528448
string GDS_START 140172
<< end >>

